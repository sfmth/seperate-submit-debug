magic
tech sky130B
magscale 1 2
timestamp 1662836958
<< obsli1 >>
rect 1104 2159 177928 178993
<< obsm1 >>
rect 1104 1708 178374 179024
<< metal2 >>
rect 662 180414 718 181214
rect 1950 180414 2006 181214
rect 3238 180414 3294 181214
rect 4526 180414 4582 181214
rect 5814 180414 5870 181214
rect 7746 180414 7802 181214
rect 9034 180414 9090 181214
rect 10322 180414 10378 181214
rect 11610 180414 11666 181214
rect 12898 180414 12954 181214
rect 14186 180414 14242 181214
rect 16118 180414 16174 181214
rect 17406 180414 17462 181214
rect 18694 180414 18750 181214
rect 19982 180414 20038 181214
rect 21270 180414 21326 181214
rect 23202 180414 23258 181214
rect 24490 180414 24546 181214
rect 25778 180414 25834 181214
rect 27066 180414 27122 181214
rect 28354 180414 28410 181214
rect 29642 180414 29698 181214
rect 31574 180414 31630 181214
rect 32862 180414 32918 181214
rect 34150 180414 34206 181214
rect 35438 180414 35494 181214
rect 36726 180414 36782 181214
rect 38014 180414 38070 181214
rect 39946 180414 40002 181214
rect 41234 180414 41290 181214
rect 42522 180414 42578 181214
rect 43810 180414 43866 181214
rect 45098 180414 45154 181214
rect 47030 180414 47086 181214
rect 48318 180414 48374 181214
rect 49606 180414 49662 181214
rect 50894 180414 50950 181214
rect 52182 180414 52238 181214
rect 53470 180414 53526 181214
rect 55402 180414 55458 181214
rect 56690 180414 56746 181214
rect 57978 180414 58034 181214
rect 59266 180414 59322 181214
rect 60554 180414 60610 181214
rect 62486 180414 62542 181214
rect 63774 180414 63830 181214
rect 65062 180414 65118 181214
rect 66350 180414 66406 181214
rect 67638 180414 67694 181214
rect 68926 180414 68982 181214
rect 70858 180414 70914 181214
rect 72146 180414 72202 181214
rect 73434 180414 73490 181214
rect 74722 180414 74778 181214
rect 76010 180414 76066 181214
rect 77942 180414 77998 181214
rect 79230 180414 79286 181214
rect 80518 180414 80574 181214
rect 81806 180414 81862 181214
rect 83094 180414 83150 181214
rect 84382 180414 84438 181214
rect 86314 180414 86370 181214
rect 87602 180414 87658 181214
rect 88890 180414 88946 181214
rect 90178 180414 90234 181214
rect 91466 180414 91522 181214
rect 93398 180414 93454 181214
rect 94686 180414 94742 181214
rect 95974 180414 96030 181214
rect 97262 180414 97318 181214
rect 98550 180414 98606 181214
rect 99838 180414 99894 181214
rect 101770 180414 101826 181214
rect 103058 180414 103114 181214
rect 104346 180414 104402 181214
rect 105634 180414 105690 181214
rect 106922 180414 106978 181214
rect 108210 180414 108266 181214
rect 110142 180414 110198 181214
rect 111430 180414 111486 181214
rect 112718 180414 112774 181214
rect 114006 180414 114062 181214
rect 115294 180414 115350 181214
rect 117226 180414 117282 181214
rect 118514 180414 118570 181214
rect 119802 180414 119858 181214
rect 121090 180414 121146 181214
rect 122378 180414 122434 181214
rect 123666 180414 123722 181214
rect 125598 180414 125654 181214
rect 126886 180414 126942 181214
rect 128174 180414 128230 181214
rect 129462 180414 129518 181214
rect 130750 180414 130806 181214
rect 132682 180414 132738 181214
rect 133970 180414 134026 181214
rect 135258 180414 135314 181214
rect 136546 180414 136602 181214
rect 137834 180414 137890 181214
rect 139122 180414 139178 181214
rect 141054 180414 141110 181214
rect 142342 180414 142398 181214
rect 143630 180414 143686 181214
rect 144918 180414 144974 181214
rect 146206 180414 146262 181214
rect 148138 180414 148194 181214
rect 149426 180414 149482 181214
rect 150714 180414 150770 181214
rect 152002 180414 152058 181214
rect 153290 180414 153346 181214
rect 154578 180414 154634 181214
rect 156510 180414 156566 181214
rect 157798 180414 157854 181214
rect 159086 180414 159142 181214
rect 160374 180414 160430 181214
rect 161662 180414 161718 181214
rect 163594 180414 163650 181214
rect 164882 180414 164938 181214
rect 166170 180414 166226 181214
rect 167458 180414 167514 181214
rect 168746 180414 168802 181214
rect 170034 180414 170090 181214
rect 171966 180414 172022 181214
rect 173254 180414 173310 181214
rect 174542 180414 174598 181214
rect 175830 180414 175886 181214
rect 177118 180414 177174 181214
rect 178406 180414 178462 181214
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 26422 0 26478 800
rect 27710 0 27766 800
rect 28998 0 29054 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 39302 0 39358 800
rect 40590 0 40646 800
rect 41878 0 41934 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 59910 0 59966 800
rect 61198 0 61254 800
rect 63130 0 63186 800
rect 64418 0 64474 800
rect 65706 0 65762 800
rect 66994 0 67050 800
rect 68282 0 68338 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72790 0 72846 800
rect 74078 0 74134 800
rect 75366 0 75422 800
rect 76654 0 76710 800
rect 78586 0 78642 800
rect 79874 0 79930 800
rect 81162 0 81218 800
rect 82450 0 82506 800
rect 83738 0 83794 800
rect 85026 0 85082 800
rect 86958 0 87014 800
rect 88246 0 88302 800
rect 89534 0 89590 800
rect 90822 0 90878 800
rect 92110 0 92166 800
rect 94042 0 94098 800
rect 95330 0 95386 800
rect 96618 0 96674 800
rect 97906 0 97962 800
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 102414 0 102470 800
rect 103702 0 103758 800
rect 104990 0 105046 800
rect 106278 0 106334 800
rect 107566 0 107622 800
rect 109498 0 109554 800
rect 110786 0 110842 800
rect 112074 0 112130 800
rect 113362 0 113418 800
rect 114650 0 114706 800
rect 115938 0 115994 800
rect 117870 0 117926 800
rect 119158 0 119214 800
rect 120446 0 120502 800
rect 121734 0 121790 800
rect 123022 0 123078 800
rect 124954 0 125010 800
rect 126242 0 126298 800
rect 127530 0 127586 800
rect 128818 0 128874 800
rect 130106 0 130162 800
rect 131394 0 131450 800
rect 133326 0 133382 800
rect 134614 0 134670 800
rect 135902 0 135958 800
rect 137190 0 137246 800
rect 138478 0 138534 800
rect 140410 0 140466 800
rect 141698 0 141754 800
rect 142986 0 143042 800
rect 144274 0 144330 800
rect 145562 0 145618 800
rect 146850 0 146906 800
rect 148782 0 148838 800
rect 150070 0 150126 800
rect 151358 0 151414 800
rect 152646 0 152702 800
rect 153934 0 153990 800
rect 155222 0 155278 800
rect 157154 0 157210 800
rect 158442 0 158498 800
rect 159730 0 159786 800
rect 161018 0 161074 800
rect 162306 0 162362 800
rect 164238 0 164294 800
rect 165526 0 165582 800
rect 166814 0 166870 800
rect 168102 0 168158 800
rect 169390 0 169446 800
rect 170678 0 170734 800
rect 172610 0 172666 800
rect 173898 0 173954 800
rect 175186 0 175242 800
rect 176474 0 176530 800
rect 177762 0 177818 800
<< obsm2 >>
rect 1308 180358 1894 180554
rect 2062 180358 3182 180554
rect 3350 180358 4470 180554
rect 4638 180358 5758 180554
rect 5926 180358 7690 180554
rect 7858 180358 8978 180554
rect 9146 180358 10266 180554
rect 10434 180358 11554 180554
rect 11722 180358 12842 180554
rect 13010 180358 14130 180554
rect 14298 180358 16062 180554
rect 16230 180358 17350 180554
rect 17518 180358 18638 180554
rect 18806 180358 19926 180554
rect 20094 180358 21214 180554
rect 21382 180358 23146 180554
rect 23314 180358 24434 180554
rect 24602 180358 25722 180554
rect 25890 180358 27010 180554
rect 27178 180358 28298 180554
rect 28466 180358 29586 180554
rect 29754 180358 31518 180554
rect 31686 180358 32806 180554
rect 32974 180358 34094 180554
rect 34262 180358 35382 180554
rect 35550 180358 36670 180554
rect 36838 180358 37958 180554
rect 38126 180358 39890 180554
rect 40058 180358 41178 180554
rect 41346 180358 42466 180554
rect 42634 180358 43754 180554
rect 43922 180358 45042 180554
rect 45210 180358 46974 180554
rect 47142 180358 48262 180554
rect 48430 180358 49550 180554
rect 49718 180358 50838 180554
rect 51006 180358 52126 180554
rect 52294 180358 53414 180554
rect 53582 180358 55346 180554
rect 55514 180358 56634 180554
rect 56802 180358 57922 180554
rect 58090 180358 59210 180554
rect 59378 180358 60498 180554
rect 60666 180358 62430 180554
rect 62598 180358 63718 180554
rect 63886 180358 65006 180554
rect 65174 180358 66294 180554
rect 66462 180358 67582 180554
rect 67750 180358 68870 180554
rect 69038 180358 70802 180554
rect 70970 180358 72090 180554
rect 72258 180358 73378 180554
rect 73546 180358 74666 180554
rect 74834 180358 75954 180554
rect 76122 180358 77886 180554
rect 78054 180358 79174 180554
rect 79342 180358 80462 180554
rect 80630 180358 81750 180554
rect 81918 180358 83038 180554
rect 83206 180358 84326 180554
rect 84494 180358 86258 180554
rect 86426 180358 87546 180554
rect 87714 180358 88834 180554
rect 89002 180358 90122 180554
rect 90290 180358 91410 180554
rect 91578 180358 93342 180554
rect 93510 180358 94630 180554
rect 94798 180358 95918 180554
rect 96086 180358 97206 180554
rect 97374 180358 98494 180554
rect 98662 180358 99782 180554
rect 99950 180358 101714 180554
rect 101882 180358 103002 180554
rect 103170 180358 104290 180554
rect 104458 180358 105578 180554
rect 105746 180358 106866 180554
rect 107034 180358 108154 180554
rect 108322 180358 110086 180554
rect 110254 180358 111374 180554
rect 111542 180358 112662 180554
rect 112830 180358 113950 180554
rect 114118 180358 115238 180554
rect 115406 180358 117170 180554
rect 117338 180358 118458 180554
rect 118626 180358 119746 180554
rect 119914 180358 121034 180554
rect 121202 180358 122322 180554
rect 122490 180358 123610 180554
rect 123778 180358 125542 180554
rect 125710 180358 126830 180554
rect 126998 180358 128118 180554
rect 128286 180358 129406 180554
rect 129574 180358 130694 180554
rect 130862 180358 132626 180554
rect 132794 180358 133914 180554
rect 134082 180358 135202 180554
rect 135370 180358 136490 180554
rect 136658 180358 137778 180554
rect 137946 180358 139066 180554
rect 139234 180358 140998 180554
rect 141166 180358 142286 180554
rect 142454 180358 143574 180554
rect 143742 180358 144862 180554
rect 145030 180358 146150 180554
rect 146318 180358 148082 180554
rect 148250 180358 149370 180554
rect 149538 180358 150658 180554
rect 150826 180358 151946 180554
rect 152114 180358 153234 180554
rect 153402 180358 154522 180554
rect 154690 180358 156454 180554
rect 156622 180358 157742 180554
rect 157910 180358 159030 180554
rect 159198 180358 160318 180554
rect 160486 180358 161606 180554
rect 161774 180358 163538 180554
rect 163706 180358 164826 180554
rect 164994 180358 166114 180554
rect 166282 180358 167402 180554
rect 167570 180358 168690 180554
rect 168858 180358 169978 180554
rect 170146 180358 171910 180554
rect 172078 180358 173198 180554
rect 173366 180358 174486 180554
rect 174654 180358 175774 180554
rect 175942 180358 177062 180554
rect 177230 180358 178350 180554
rect 1308 856 178406 180358
rect 1418 734 2538 856
rect 2706 734 3826 856
rect 3994 734 5114 856
rect 5282 734 6402 856
rect 6570 734 8334 856
rect 8502 734 9622 856
rect 9790 734 10910 856
rect 11078 734 12198 856
rect 12366 734 13486 856
rect 13654 734 14774 856
rect 14942 734 16706 856
rect 16874 734 17994 856
rect 18162 734 19282 856
rect 19450 734 20570 856
rect 20738 734 21858 856
rect 22026 734 23790 856
rect 23958 734 25078 856
rect 25246 734 26366 856
rect 26534 734 27654 856
rect 27822 734 28942 856
rect 29110 734 30230 856
rect 30398 734 32162 856
rect 32330 734 33450 856
rect 33618 734 34738 856
rect 34906 734 36026 856
rect 36194 734 37314 856
rect 37482 734 39246 856
rect 39414 734 40534 856
rect 40702 734 41822 856
rect 41990 734 43110 856
rect 43278 734 44398 856
rect 44566 734 45686 856
rect 45854 734 47618 856
rect 47786 734 48906 856
rect 49074 734 50194 856
rect 50362 734 51482 856
rect 51650 734 52770 856
rect 52938 734 54702 856
rect 54870 734 55990 856
rect 56158 734 57278 856
rect 57446 734 58566 856
rect 58734 734 59854 856
rect 60022 734 61142 856
rect 61310 734 63074 856
rect 63242 734 64362 856
rect 64530 734 65650 856
rect 65818 734 66938 856
rect 67106 734 68226 856
rect 68394 734 70158 856
rect 70326 734 71446 856
rect 71614 734 72734 856
rect 72902 734 74022 856
rect 74190 734 75310 856
rect 75478 734 76598 856
rect 76766 734 78530 856
rect 78698 734 79818 856
rect 79986 734 81106 856
rect 81274 734 82394 856
rect 82562 734 83682 856
rect 83850 734 84970 856
rect 85138 734 86902 856
rect 87070 734 88190 856
rect 88358 734 89478 856
rect 89646 734 90766 856
rect 90934 734 92054 856
rect 92222 734 93986 856
rect 94154 734 95274 856
rect 95442 734 96562 856
rect 96730 734 97850 856
rect 98018 734 99138 856
rect 99306 734 100426 856
rect 100594 734 102358 856
rect 102526 734 103646 856
rect 103814 734 104934 856
rect 105102 734 106222 856
rect 106390 734 107510 856
rect 107678 734 109442 856
rect 109610 734 110730 856
rect 110898 734 112018 856
rect 112186 734 113306 856
rect 113474 734 114594 856
rect 114762 734 115882 856
rect 116050 734 117814 856
rect 117982 734 119102 856
rect 119270 734 120390 856
rect 120558 734 121678 856
rect 121846 734 122966 856
rect 123134 734 124898 856
rect 125066 734 126186 856
rect 126354 734 127474 856
rect 127642 734 128762 856
rect 128930 734 130050 856
rect 130218 734 131338 856
rect 131506 734 133270 856
rect 133438 734 134558 856
rect 134726 734 135846 856
rect 136014 734 137134 856
rect 137302 734 138422 856
rect 138590 734 140354 856
rect 140522 734 141642 856
rect 141810 734 142930 856
rect 143098 734 144218 856
rect 144386 734 145506 856
rect 145674 734 146794 856
rect 146962 734 148726 856
rect 148894 734 150014 856
rect 150182 734 151302 856
rect 151470 734 152590 856
rect 152758 734 153878 856
rect 154046 734 155166 856
rect 155334 734 157098 856
rect 157266 734 158386 856
rect 158554 734 159674 856
rect 159842 734 160962 856
rect 161130 734 162250 856
rect 162418 734 164182 856
rect 164350 734 165470 856
rect 165638 734 166758 856
rect 166926 734 168046 856
rect 168214 734 169334 856
rect 169502 734 170622 856
rect 170790 734 172554 856
rect 172722 734 173842 856
rect 174010 734 175130 856
rect 175298 734 176418 856
rect 176586 734 177706 856
rect 177874 734 178406 856
<< metal3 >>
rect 0 180208 800 180328
rect 178270 179528 179070 179648
rect 0 178848 800 178968
rect 178270 178168 179070 178288
rect 0 177488 800 177608
rect 178270 176808 179070 176928
rect 0 176128 800 176248
rect 178270 175448 179070 175568
rect 0 174768 800 174888
rect 178270 174088 179070 174208
rect 0 173408 800 173528
rect 178270 172048 179070 172168
rect 0 171368 800 171488
rect 178270 170688 179070 170808
rect 0 170008 800 170128
rect 178270 169328 179070 169448
rect 0 168648 800 168768
rect 178270 167968 179070 168088
rect 0 167288 800 167408
rect 178270 166608 179070 166728
rect 0 165928 800 166048
rect 178270 165248 179070 165368
rect 0 163888 800 164008
rect 178270 163208 179070 163328
rect 0 162528 800 162648
rect 178270 161848 179070 161968
rect 0 161168 800 161288
rect 178270 160488 179070 160608
rect 0 159808 800 159928
rect 178270 159128 179070 159248
rect 0 158448 800 158568
rect 178270 157768 179070 157888
rect 0 157088 800 157208
rect 178270 155728 179070 155848
rect 0 155048 800 155168
rect 178270 154368 179070 154488
rect 0 153688 800 153808
rect 178270 153008 179070 153128
rect 0 152328 800 152448
rect 178270 151648 179070 151768
rect 0 150968 800 151088
rect 178270 150288 179070 150408
rect 0 149608 800 149728
rect 178270 148928 179070 149048
rect 0 147568 800 147688
rect 178270 146888 179070 147008
rect 0 146208 800 146328
rect 178270 145528 179070 145648
rect 0 144848 800 144968
rect 178270 144168 179070 144288
rect 0 143488 800 143608
rect 178270 142808 179070 142928
rect 0 142128 800 142248
rect 178270 141448 179070 141568
rect 0 140768 800 140888
rect 178270 139408 179070 139528
rect 0 138728 800 138848
rect 178270 138048 179070 138168
rect 0 137368 800 137488
rect 178270 136688 179070 136808
rect 0 136008 800 136128
rect 178270 135328 179070 135448
rect 0 134648 800 134768
rect 178270 133968 179070 134088
rect 0 133288 800 133408
rect 178270 132608 179070 132728
rect 0 131928 800 132048
rect 178270 130568 179070 130688
rect 0 129888 800 130008
rect 178270 129208 179070 129328
rect 0 128528 800 128648
rect 178270 127848 179070 127968
rect 0 127168 800 127288
rect 178270 126488 179070 126608
rect 0 125808 800 125928
rect 178270 125128 179070 125248
rect 0 124448 800 124568
rect 178270 123088 179070 123208
rect 0 122408 800 122528
rect 178270 121728 179070 121848
rect 0 121048 800 121168
rect 178270 120368 179070 120488
rect 0 119688 800 119808
rect 178270 119008 179070 119128
rect 0 118328 800 118448
rect 178270 117648 179070 117768
rect 0 116968 800 117088
rect 178270 116288 179070 116408
rect 0 115608 800 115728
rect 178270 114248 179070 114368
rect 0 113568 800 113688
rect 178270 112888 179070 113008
rect 0 112208 800 112328
rect 178270 111528 179070 111648
rect 0 110848 800 110968
rect 178270 110168 179070 110288
rect 0 109488 800 109608
rect 178270 108808 179070 108928
rect 0 108128 800 108248
rect 178270 107448 179070 107568
rect 0 106088 800 106208
rect 178270 105408 179070 105528
rect 0 104728 800 104848
rect 178270 104048 179070 104168
rect 0 103368 800 103488
rect 178270 102688 179070 102808
rect 0 102008 800 102128
rect 178270 101328 179070 101448
rect 0 100648 800 100768
rect 178270 99968 179070 100088
rect 0 99288 800 99408
rect 178270 97928 179070 98048
rect 0 97248 800 97368
rect 178270 96568 179070 96688
rect 0 95888 800 96008
rect 178270 95208 179070 95328
rect 0 94528 800 94648
rect 178270 93848 179070 93968
rect 0 93168 800 93288
rect 178270 92488 179070 92608
rect 0 91808 800 91928
rect 178270 91128 179070 91248
rect 0 89768 800 89888
rect 178270 89088 179070 89208
rect 0 88408 800 88528
rect 178270 87728 179070 87848
rect 0 87048 800 87168
rect 178270 86368 179070 86488
rect 0 85688 800 85808
rect 178270 85008 179070 85128
rect 0 84328 800 84448
rect 178270 83648 179070 83768
rect 0 82968 800 83088
rect 178270 81608 179070 81728
rect 0 80928 800 81048
rect 178270 80248 179070 80368
rect 0 79568 800 79688
rect 178270 78888 179070 79008
rect 0 78208 800 78328
rect 178270 77528 179070 77648
rect 0 76848 800 76968
rect 178270 76168 179070 76288
rect 0 75488 800 75608
rect 178270 74808 179070 74928
rect 0 73448 800 73568
rect 178270 72768 179070 72888
rect 0 72088 800 72208
rect 178270 71408 179070 71528
rect 0 70728 800 70848
rect 178270 70048 179070 70168
rect 0 69368 800 69488
rect 178270 68688 179070 68808
rect 0 68008 800 68128
rect 178270 67328 179070 67448
rect 0 66648 800 66768
rect 178270 65288 179070 65408
rect 0 64608 800 64728
rect 178270 63928 179070 64048
rect 0 63248 800 63368
rect 178270 62568 179070 62688
rect 0 61888 800 62008
rect 178270 61208 179070 61328
rect 0 60528 800 60648
rect 178270 59848 179070 59968
rect 0 59168 800 59288
rect 178270 58488 179070 58608
rect 0 57808 800 57928
rect 178270 56448 179070 56568
rect 0 55768 800 55888
rect 178270 55088 179070 55208
rect 0 54408 800 54528
rect 178270 53728 179070 53848
rect 0 53048 800 53168
rect 178270 52368 179070 52488
rect 0 51688 800 51808
rect 178270 51008 179070 51128
rect 0 50328 800 50448
rect 178270 48968 179070 49088
rect 0 48288 800 48408
rect 178270 47608 179070 47728
rect 0 46928 800 47048
rect 178270 46248 179070 46368
rect 0 45568 800 45688
rect 178270 44888 179070 45008
rect 0 44208 800 44328
rect 178270 43528 179070 43648
rect 0 42848 800 42968
rect 178270 42168 179070 42288
rect 0 41488 800 41608
rect 178270 40128 179070 40248
rect 0 39448 800 39568
rect 178270 38768 179070 38888
rect 0 38088 800 38208
rect 178270 37408 179070 37528
rect 0 36728 800 36848
rect 178270 36048 179070 36168
rect 0 35368 800 35488
rect 178270 34688 179070 34808
rect 0 34008 800 34128
rect 178270 33328 179070 33448
rect 0 31968 800 32088
rect 178270 31288 179070 31408
rect 0 30608 800 30728
rect 178270 29928 179070 30048
rect 0 29248 800 29368
rect 178270 28568 179070 28688
rect 0 27888 800 28008
rect 178270 27208 179070 27328
rect 0 26528 800 26648
rect 178270 25848 179070 25968
rect 0 25168 800 25288
rect 178270 23808 179070 23928
rect 0 23128 800 23248
rect 178270 22448 179070 22568
rect 0 21768 800 21888
rect 178270 21088 179070 21208
rect 0 20408 800 20528
rect 178270 19728 179070 19848
rect 0 19048 800 19168
rect 178270 18368 179070 18488
rect 0 17688 800 17808
rect 178270 17008 179070 17128
rect 0 15648 800 15768
rect 178270 14968 179070 15088
rect 0 14288 800 14408
rect 178270 13608 179070 13728
rect 0 12928 800 13048
rect 178270 12248 179070 12368
rect 0 11568 800 11688
rect 178270 10888 179070 11008
rect 0 10208 800 10328
rect 178270 9528 179070 9648
rect 0 8848 800 8968
rect 178270 7488 179070 7608
rect 0 6808 800 6928
rect 178270 6128 179070 6248
rect 0 5448 800 5568
rect 178270 4768 179070 4888
rect 0 4088 800 4208
rect 178270 3408 179070 3528
rect 0 2728 800 2848
rect 178270 2048 179070 2168
rect 0 1368 800 1488
rect 178270 688 179070 808
<< obsm3 >>
rect 800 179448 178190 179621
rect 800 179048 178270 179448
rect 880 178768 178270 179048
rect 800 178368 178270 178768
rect 800 178088 178190 178368
rect 800 177688 178270 178088
rect 880 177408 178270 177688
rect 800 177008 178270 177408
rect 800 176728 178190 177008
rect 800 176328 178270 176728
rect 880 176048 178270 176328
rect 800 175648 178270 176048
rect 800 175368 178190 175648
rect 800 174968 178270 175368
rect 880 174688 178270 174968
rect 800 174288 178270 174688
rect 800 174008 178190 174288
rect 800 173608 178270 174008
rect 880 173328 178270 173608
rect 800 172248 178270 173328
rect 800 171968 178190 172248
rect 800 171568 178270 171968
rect 880 171288 178270 171568
rect 800 170888 178270 171288
rect 800 170608 178190 170888
rect 800 170208 178270 170608
rect 880 169928 178270 170208
rect 800 169528 178270 169928
rect 800 169248 178190 169528
rect 800 168848 178270 169248
rect 880 168568 178270 168848
rect 800 168168 178270 168568
rect 800 167888 178190 168168
rect 800 167488 178270 167888
rect 880 167208 178270 167488
rect 800 166808 178270 167208
rect 800 166528 178190 166808
rect 800 166128 178270 166528
rect 880 165848 178270 166128
rect 800 165448 178270 165848
rect 800 165168 178190 165448
rect 800 164088 178270 165168
rect 880 163808 178270 164088
rect 800 163408 178270 163808
rect 800 163128 178190 163408
rect 800 162728 178270 163128
rect 880 162448 178270 162728
rect 800 162048 178270 162448
rect 800 161768 178190 162048
rect 800 161368 178270 161768
rect 880 161088 178270 161368
rect 800 160688 178270 161088
rect 800 160408 178190 160688
rect 800 160008 178270 160408
rect 880 159728 178270 160008
rect 800 159328 178270 159728
rect 800 159048 178190 159328
rect 800 158648 178270 159048
rect 880 158368 178270 158648
rect 800 157968 178270 158368
rect 800 157688 178190 157968
rect 800 157288 178270 157688
rect 880 157008 178270 157288
rect 800 155928 178270 157008
rect 800 155648 178190 155928
rect 800 155248 178270 155648
rect 880 154968 178270 155248
rect 800 154568 178270 154968
rect 800 154288 178190 154568
rect 800 153888 178270 154288
rect 880 153608 178270 153888
rect 800 153208 178270 153608
rect 800 152928 178190 153208
rect 800 152528 178270 152928
rect 880 152248 178270 152528
rect 800 151848 178270 152248
rect 800 151568 178190 151848
rect 800 151168 178270 151568
rect 880 150888 178270 151168
rect 800 150488 178270 150888
rect 800 150208 178190 150488
rect 800 149808 178270 150208
rect 880 149528 178270 149808
rect 800 149128 178270 149528
rect 800 148848 178190 149128
rect 800 147768 178270 148848
rect 880 147488 178270 147768
rect 800 147088 178270 147488
rect 800 146808 178190 147088
rect 800 146408 178270 146808
rect 880 146128 178270 146408
rect 800 145728 178270 146128
rect 800 145448 178190 145728
rect 800 145048 178270 145448
rect 880 144768 178270 145048
rect 800 144368 178270 144768
rect 800 144088 178190 144368
rect 800 143688 178270 144088
rect 880 143408 178270 143688
rect 800 143008 178270 143408
rect 800 142728 178190 143008
rect 800 142328 178270 142728
rect 880 142048 178270 142328
rect 800 141648 178270 142048
rect 800 141368 178190 141648
rect 800 140968 178270 141368
rect 880 140688 178270 140968
rect 800 139608 178270 140688
rect 800 139328 178190 139608
rect 800 138928 178270 139328
rect 880 138648 178270 138928
rect 800 138248 178270 138648
rect 800 137968 178190 138248
rect 800 137568 178270 137968
rect 880 137288 178270 137568
rect 800 136888 178270 137288
rect 800 136608 178190 136888
rect 800 136208 178270 136608
rect 880 135928 178270 136208
rect 800 135528 178270 135928
rect 800 135248 178190 135528
rect 800 134848 178270 135248
rect 880 134568 178270 134848
rect 800 134168 178270 134568
rect 800 133888 178190 134168
rect 800 133488 178270 133888
rect 880 133208 178270 133488
rect 800 132808 178270 133208
rect 800 132528 178190 132808
rect 800 132128 178270 132528
rect 880 131848 178270 132128
rect 800 130768 178270 131848
rect 800 130488 178190 130768
rect 800 130088 178270 130488
rect 880 129808 178270 130088
rect 800 129408 178270 129808
rect 800 129128 178190 129408
rect 800 128728 178270 129128
rect 880 128448 178270 128728
rect 800 128048 178270 128448
rect 800 127768 178190 128048
rect 800 127368 178270 127768
rect 880 127088 178270 127368
rect 800 126688 178270 127088
rect 800 126408 178190 126688
rect 800 126008 178270 126408
rect 880 125728 178270 126008
rect 800 125328 178270 125728
rect 800 125048 178190 125328
rect 800 124648 178270 125048
rect 880 124368 178270 124648
rect 800 123288 178270 124368
rect 800 123008 178190 123288
rect 800 122608 178270 123008
rect 880 122328 178270 122608
rect 800 121928 178270 122328
rect 800 121648 178190 121928
rect 800 121248 178270 121648
rect 880 120968 178270 121248
rect 800 120568 178270 120968
rect 800 120288 178190 120568
rect 800 119888 178270 120288
rect 880 119608 178270 119888
rect 800 119208 178270 119608
rect 800 118928 178190 119208
rect 800 118528 178270 118928
rect 880 118248 178270 118528
rect 800 117848 178270 118248
rect 800 117568 178190 117848
rect 800 117168 178270 117568
rect 880 116888 178270 117168
rect 800 116488 178270 116888
rect 800 116208 178190 116488
rect 800 115808 178270 116208
rect 880 115528 178270 115808
rect 800 114448 178270 115528
rect 800 114168 178190 114448
rect 800 113768 178270 114168
rect 880 113488 178270 113768
rect 800 113088 178270 113488
rect 800 112808 178190 113088
rect 800 112408 178270 112808
rect 880 112128 178270 112408
rect 800 111728 178270 112128
rect 800 111448 178190 111728
rect 800 111048 178270 111448
rect 880 110768 178270 111048
rect 800 110368 178270 110768
rect 800 110088 178190 110368
rect 800 109688 178270 110088
rect 880 109408 178270 109688
rect 800 109008 178270 109408
rect 800 108728 178190 109008
rect 800 108328 178270 108728
rect 880 108048 178270 108328
rect 800 107648 178270 108048
rect 800 107368 178190 107648
rect 800 106288 178270 107368
rect 880 106008 178270 106288
rect 800 105608 178270 106008
rect 800 105328 178190 105608
rect 800 104928 178270 105328
rect 880 104648 178270 104928
rect 800 104248 178270 104648
rect 800 103968 178190 104248
rect 800 103568 178270 103968
rect 880 103288 178270 103568
rect 800 102888 178270 103288
rect 800 102608 178190 102888
rect 800 102208 178270 102608
rect 880 101928 178270 102208
rect 800 101528 178270 101928
rect 800 101248 178190 101528
rect 800 100848 178270 101248
rect 880 100568 178270 100848
rect 800 100168 178270 100568
rect 800 99888 178190 100168
rect 800 99488 178270 99888
rect 880 99208 178270 99488
rect 800 98128 178270 99208
rect 800 97848 178190 98128
rect 800 97448 178270 97848
rect 880 97168 178270 97448
rect 800 96768 178270 97168
rect 800 96488 178190 96768
rect 800 96088 178270 96488
rect 880 95808 178270 96088
rect 800 95408 178270 95808
rect 800 95128 178190 95408
rect 800 94728 178270 95128
rect 880 94448 178270 94728
rect 800 94048 178270 94448
rect 800 93768 178190 94048
rect 800 93368 178270 93768
rect 880 93088 178270 93368
rect 800 92688 178270 93088
rect 800 92408 178190 92688
rect 800 92008 178270 92408
rect 880 91728 178270 92008
rect 800 91328 178270 91728
rect 800 91048 178190 91328
rect 800 89968 178270 91048
rect 880 89688 178270 89968
rect 800 89288 178270 89688
rect 800 89008 178190 89288
rect 800 88608 178270 89008
rect 880 88328 178270 88608
rect 800 87928 178270 88328
rect 800 87648 178190 87928
rect 800 87248 178270 87648
rect 880 86968 178270 87248
rect 800 86568 178270 86968
rect 800 86288 178190 86568
rect 800 85888 178270 86288
rect 880 85608 178270 85888
rect 800 85208 178270 85608
rect 800 84928 178190 85208
rect 800 84528 178270 84928
rect 880 84248 178270 84528
rect 800 83848 178270 84248
rect 800 83568 178190 83848
rect 800 83168 178270 83568
rect 880 82888 178270 83168
rect 800 81808 178270 82888
rect 800 81528 178190 81808
rect 800 81128 178270 81528
rect 880 80848 178270 81128
rect 800 80448 178270 80848
rect 800 80168 178190 80448
rect 800 79768 178270 80168
rect 880 79488 178270 79768
rect 800 79088 178270 79488
rect 800 78808 178190 79088
rect 800 78408 178270 78808
rect 880 78128 178270 78408
rect 800 77728 178270 78128
rect 800 77448 178190 77728
rect 800 77048 178270 77448
rect 880 76768 178270 77048
rect 800 76368 178270 76768
rect 800 76088 178190 76368
rect 800 75688 178270 76088
rect 880 75408 178270 75688
rect 800 75008 178270 75408
rect 800 74728 178190 75008
rect 800 73648 178270 74728
rect 880 73368 178270 73648
rect 800 72968 178270 73368
rect 800 72688 178190 72968
rect 800 72288 178270 72688
rect 880 72008 178270 72288
rect 800 71608 178270 72008
rect 800 71328 178190 71608
rect 800 70928 178270 71328
rect 880 70648 178270 70928
rect 800 70248 178270 70648
rect 800 69968 178190 70248
rect 800 69568 178270 69968
rect 880 69288 178270 69568
rect 800 68888 178270 69288
rect 800 68608 178190 68888
rect 800 68208 178270 68608
rect 880 67928 178270 68208
rect 800 67528 178270 67928
rect 800 67248 178190 67528
rect 800 66848 178270 67248
rect 880 66568 178270 66848
rect 800 65488 178270 66568
rect 800 65208 178190 65488
rect 800 64808 178270 65208
rect 880 64528 178270 64808
rect 800 64128 178270 64528
rect 800 63848 178190 64128
rect 800 63448 178270 63848
rect 880 63168 178270 63448
rect 800 62768 178270 63168
rect 800 62488 178190 62768
rect 800 62088 178270 62488
rect 880 61808 178270 62088
rect 800 61408 178270 61808
rect 800 61128 178190 61408
rect 800 60728 178270 61128
rect 880 60448 178270 60728
rect 800 60048 178270 60448
rect 800 59768 178190 60048
rect 800 59368 178270 59768
rect 880 59088 178270 59368
rect 800 58688 178270 59088
rect 800 58408 178190 58688
rect 800 58008 178270 58408
rect 880 57728 178270 58008
rect 800 56648 178270 57728
rect 800 56368 178190 56648
rect 800 55968 178270 56368
rect 880 55688 178270 55968
rect 800 55288 178270 55688
rect 800 55008 178190 55288
rect 800 54608 178270 55008
rect 880 54328 178270 54608
rect 800 53928 178270 54328
rect 800 53648 178190 53928
rect 800 53248 178270 53648
rect 880 52968 178270 53248
rect 800 52568 178270 52968
rect 800 52288 178190 52568
rect 800 51888 178270 52288
rect 880 51608 178270 51888
rect 800 51208 178270 51608
rect 800 50928 178190 51208
rect 800 50528 178270 50928
rect 880 50248 178270 50528
rect 800 49168 178270 50248
rect 800 48888 178190 49168
rect 800 48488 178270 48888
rect 880 48208 178270 48488
rect 800 47808 178270 48208
rect 800 47528 178190 47808
rect 800 47128 178270 47528
rect 880 46848 178270 47128
rect 800 46448 178270 46848
rect 800 46168 178190 46448
rect 800 45768 178270 46168
rect 880 45488 178270 45768
rect 800 45088 178270 45488
rect 800 44808 178190 45088
rect 800 44408 178270 44808
rect 880 44128 178270 44408
rect 800 43728 178270 44128
rect 800 43448 178190 43728
rect 800 43048 178270 43448
rect 880 42768 178270 43048
rect 800 42368 178270 42768
rect 800 42088 178190 42368
rect 800 41688 178270 42088
rect 880 41408 178270 41688
rect 800 40328 178270 41408
rect 800 40048 178190 40328
rect 800 39648 178270 40048
rect 880 39368 178270 39648
rect 800 38968 178270 39368
rect 800 38688 178190 38968
rect 800 38288 178270 38688
rect 880 38008 178270 38288
rect 800 37608 178270 38008
rect 800 37328 178190 37608
rect 800 36928 178270 37328
rect 880 36648 178270 36928
rect 800 36248 178270 36648
rect 800 35968 178190 36248
rect 800 35568 178270 35968
rect 880 35288 178270 35568
rect 800 34888 178270 35288
rect 800 34608 178190 34888
rect 800 34208 178270 34608
rect 880 33928 178270 34208
rect 800 33528 178270 33928
rect 800 33248 178190 33528
rect 800 32168 178270 33248
rect 880 31888 178270 32168
rect 800 31488 178270 31888
rect 800 31208 178190 31488
rect 800 30808 178270 31208
rect 880 30528 178270 30808
rect 800 30128 178270 30528
rect 800 29848 178190 30128
rect 800 29448 178270 29848
rect 880 29168 178270 29448
rect 800 28768 178270 29168
rect 800 28488 178190 28768
rect 800 28088 178270 28488
rect 880 27808 178270 28088
rect 800 27408 178270 27808
rect 800 27128 178190 27408
rect 800 26728 178270 27128
rect 880 26448 178270 26728
rect 800 26048 178270 26448
rect 800 25768 178190 26048
rect 800 25368 178270 25768
rect 880 25088 178270 25368
rect 800 24008 178270 25088
rect 800 23728 178190 24008
rect 800 23328 178270 23728
rect 880 23048 178270 23328
rect 800 22648 178270 23048
rect 800 22368 178190 22648
rect 800 21968 178270 22368
rect 880 21688 178270 21968
rect 800 21288 178270 21688
rect 800 21008 178190 21288
rect 800 20608 178270 21008
rect 880 20328 178270 20608
rect 800 19928 178270 20328
rect 800 19648 178190 19928
rect 800 19248 178270 19648
rect 880 18968 178270 19248
rect 800 18568 178270 18968
rect 800 18288 178190 18568
rect 800 17888 178270 18288
rect 880 17608 178270 17888
rect 800 17208 178270 17608
rect 800 16928 178190 17208
rect 800 15848 178270 16928
rect 880 15568 178270 15848
rect 800 15168 178270 15568
rect 800 14888 178190 15168
rect 800 14488 178270 14888
rect 880 14208 178270 14488
rect 800 13808 178270 14208
rect 800 13528 178190 13808
rect 800 13128 178270 13528
rect 880 12848 178270 13128
rect 800 12448 178270 12848
rect 800 12168 178190 12448
rect 800 11768 178270 12168
rect 880 11488 178270 11768
rect 800 11088 178270 11488
rect 800 10808 178190 11088
rect 800 10408 178270 10808
rect 880 10128 178270 10408
rect 800 9728 178270 10128
rect 800 9448 178190 9728
rect 800 9048 178270 9448
rect 880 8768 178270 9048
rect 800 7688 178270 8768
rect 800 7408 178190 7688
rect 800 7008 178270 7408
rect 880 6728 178270 7008
rect 800 6328 178270 6728
rect 800 6048 178190 6328
rect 800 5648 178270 6048
rect 880 5368 178270 5648
rect 800 4968 178270 5368
rect 800 4688 178190 4968
rect 800 4288 178270 4688
rect 880 4008 178270 4288
rect 800 3608 178270 4008
rect 800 3328 178190 3608
rect 800 2928 178270 3328
rect 880 2648 178270 2928
rect 800 2248 178270 2648
rect 800 1968 178190 2248
rect 800 1568 178270 1968
rect 880 1395 178270 1568
<< metal4 >>
rect 4208 2128 4528 179024
rect 19568 2128 19888 179024
rect 34928 2128 35248 179024
rect 50288 2128 50608 179024
rect 65648 2128 65968 179024
rect 81008 2128 81328 179024
rect 96368 2128 96688 179024
rect 111728 2128 112048 179024
rect 127088 2128 127408 179024
rect 142448 2128 142768 179024
rect 157808 2128 158128 179024
rect 173168 2128 173488 179024
<< obsm4 >>
rect 5579 8875 19488 177037
rect 19968 8875 34848 177037
rect 35328 8875 50208 177037
rect 50688 8875 65568 177037
rect 66048 8875 80928 177037
rect 81408 8875 96288 177037
rect 96768 8875 111648 177037
rect 112128 8875 127008 177037
rect 127488 8875 142368 177037
rect 142848 8875 157728 177037
rect 158208 8875 164069 177037
<< labels >>
rlabel metal3 s 178270 76168 179070 76288 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 68926 180414 68982 181214 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 148138 180414 148194 181214 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 178270 83648 179070 83768 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 178270 132608 179070 132728 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 169390 0 169446 800 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 178270 43528 179070 43648 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 162306 0 162362 800 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 119802 180414 119858 181214 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 136546 180414 136602 181214 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 110142 180414 110198 181214 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 41234 180414 41290 181214 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 io_in[22]
port 15 nsew signal input
rlabel metal3 s 178270 2048 179070 2168 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 32862 180414 32918 181214 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 178270 175448 179070 175568 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 178270 93848 179070 93968 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 10322 180414 10378 181214 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 161168 800 161288 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 105634 180414 105690 181214 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 178270 77528 179070 77648 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 178270 33328 179070 33448 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 178270 80248 179070 80368 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 166170 180414 166226 181214 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 178270 52368 179070 52488 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 178270 10888 179070 11008 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 23202 180414 23258 181214 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 178270 125128 179070 125248 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 0 173408 800 173528 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 53470 180414 53526 181214 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 146206 180414 146262 181214 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 io_oeb[14]
port 44 nsew signal output
rlabel metal3 s 178270 72768 179070 72888 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 178270 27208 179070 27328 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 178406 180414 178462 181214 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 178270 97928 179070 98048 6 io_oeb[18]
port 48 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 0 144848 800 144968 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 io_oeb[20]
port 51 nsew signal output
rlabel metal3 s 178270 95208 179070 95328 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 123022 0 123078 800 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 0 134648 800 134768 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 174542 180414 174598 181214 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 21270 180414 21326 181214 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 159086 180414 159142 181214 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 124448 800 124568 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 88890 180414 88946 181214 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 178270 14968 179070 15088 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 178270 23808 179070 23928 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 178270 61208 179070 61328 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 3238 180414 3294 181214 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 178270 46248 179070 46368 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 178270 22448 179070 22568 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 142342 180414 142398 181214 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 14186 180414 14242 181214 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 0 163888 800 164008 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 121090 180414 121146 181214 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 178270 4768 179070 4888 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 0 177488 800 177608 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 70858 180414 70914 181214 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 177118 180414 177174 181214 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 49606 180414 49662 181214 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 103058 180414 103114 181214 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 36726 180414 36782 181214 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 178270 47608 179070 47728 6 io_out[22]
port 91 nsew signal output
rlabel metal3 s 178270 119008 179070 119128 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 178270 13608 179070 13728 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 38014 180414 38070 181214 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 178270 163208 179070 163328 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 178270 40128 179070 40248 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 110848 800 110968 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 178270 105408 179070 105528 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 74722 180414 74778 181214 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 178270 29928 179070 30048 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 178270 142808 179070 142928 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 178270 151648 179070 151768 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 0 174768 800 174888 6 la_data_in[0]
port 115 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 la_data_in[100]
port 116 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_data_in[101]
port 117 nsew signal input
rlabel metal3 s 178270 92488 179070 92608 6 la_data_in[102]
port 118 nsew signal input
rlabel metal3 s 178270 160488 179070 160608 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 101770 180414 101826 181214 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 106922 180414 106978 181214 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal3 s 178270 126488 179070 126608 6 la_data_in[109]
port 125 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 la_data_in[10]
port 126 nsew signal input
rlabel metal3 s 0 176128 800 176248 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 29642 180414 29698 181214 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal3 s 178270 127848 179070 127968 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 52182 180414 52238 181214 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 128174 180414 128230 181214 6 la_data_in[119]
port 136 nsew signal input
rlabel metal3 s 178270 99968 179070 100088 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 144918 180414 144974 181214 6 la_data_in[120]
port 138 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 la_data_in[121]
port 139 nsew signal input
rlabel metal3 s 178270 102688 179070 102808 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 98550 180414 98606 181214 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 166814 0 166870 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 la_data_in[126]
port 144 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[127]
port 145 nsew signal input
rlabel metal3 s 178270 108808 179070 108928 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 133970 180414 134026 181214 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 662 180414 718 181214 6 la_data_in[14]
port 148 nsew signal input
rlabel metal3 s 178270 18368 179070 18488 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal3 s 178270 139408 179070 139528 6 la_data_in[17]
port 151 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 la_data_in[18]
port 152 nsew signal input
rlabel metal3 s 178270 58488 179070 58608 6 la_data_in[19]
port 153 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal3 s 178270 155728 179070 155848 6 la_data_in[21]
port 156 nsew signal input
rlabel metal3 s 178270 70048 179070 70168 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 16118 180414 16174 181214 6 la_data_in[25]
port 160 nsew signal input
rlabel metal3 s 178270 161848 179070 161968 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal3 s 178270 17008 179070 17128 6 la_data_in[28]
port 163 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 45098 180414 45154 181214 6 la_data_in[33]
port 169 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_data_in[34]
port 170 nsew signal input
rlabel metal3 s 178270 12248 179070 12368 6 la_data_in[35]
port 171 nsew signal input
rlabel metal3 s 178270 86368 179070 86488 6 la_data_in[36]
port 172 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_data_in[37]
port 173 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 11610 180414 11666 181214 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 59266 180414 59322 181214 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 55402 180414 55458 181214 6 la_data_in[40]
port 177 nsew signal input
rlabel metal3 s 178270 89088 179070 89208 6 la_data_in[41]
port 178 nsew signal input
rlabel metal3 s 178270 112888 179070 113008 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal3 s 178270 25848 179070 25968 6 la_data_in[44]
port 181 nsew signal input
rlabel metal3 s 178270 6128 179070 6248 6 la_data_in[45]
port 182 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 175830 180414 175886 181214 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 163594 180414 163650 181214 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal3 s 178270 104048 179070 104168 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 112718 180414 112774 181214 6 la_data_in[54]
port 192 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 131394 0 131450 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal3 s 178270 114248 179070 114368 6 la_data_in[57]
port 195 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 la_data_in[58]
port 196 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 73434 180414 73490 181214 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 77942 180414 77998 181214 6 la_data_in[61]
port 200 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 4526 180414 4582 181214 6 la_data_in[63]
port 202 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 la_data_in[64]
port 203 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 164882 180414 164938 181214 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 65062 180414 65118 181214 6 la_data_in[67]
port 206 nsew signal input
rlabel metal3 s 178270 176808 179070 176928 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 84382 180414 84438 181214 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 104346 180414 104402 181214 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 56690 180414 56746 181214 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 108210 180414 108266 181214 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 167458 180414 167514 181214 6 la_data_in[73]
port 213 nsew signal input
rlabel metal3 s 0 180208 800 180328 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 83094 180414 83150 181214 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 67638 180414 67694 181214 6 la_data_in[76]
port 216 nsew signal input
rlabel metal3 s 0 150968 800 151088 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 173254 180414 173310 181214 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 75366 0 75422 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal3 s 178270 174088 179070 174208 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 161662 180414 161718 181214 6 la_data_in[80]
port 221 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 la_data_in[81]
port 222 nsew signal input
rlabel metal3 s 0 125808 800 125928 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 39946 180414 40002 181214 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal3 s 178270 44888 179070 45008 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 176474 0 176530 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 76010 180414 76066 181214 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 la_data_in[89]
port 230 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 99838 180414 99894 181214 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 94686 180414 94742 181214 6 la_data_in[92]
port 234 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 150714 180414 150770 181214 6 la_data_in[94]
port 236 nsew signal input
rlabel metal3 s 178270 53728 179070 53848 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 la_data_in[98]
port 240 nsew signal input
rlabel metal3 s 178270 688 179070 808 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 63774 180414 63830 181214 6 la_data_in[9]
port 242 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 31574 180414 31630 181214 6 la_data_out[100]
port 244 nsew signal output
rlabel metal3 s 0 146208 800 146328 6 la_data_out[101]
port 245 nsew signal output
rlabel metal3 s 0 140768 800 140888 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 121734 0 121790 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal3 s 178270 110168 179070 110288 6 la_data_out[104]
port 248 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 la_data_out[105]
port 249 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 la_data_out[106]
port 250 nsew signal output
rlabel metal3 s 178270 51008 179070 51128 6 la_data_out[107]
port 251 nsew signal output
rlabel metal3 s 0 162528 800 162648 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 168746 180414 168802 181214 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 137834 180414 137890 181214 6 la_data_out[111]
port 256 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 la_data_out[112]
port 257 nsew signal output
rlabel metal3 s 178270 153008 179070 153128 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 60554 180414 60610 181214 6 la_data_out[114]
port 259 nsew signal output
rlabel metal3 s 178270 120368 179070 120488 6 la_data_out[115]
port 260 nsew signal output
rlabel metal3 s 0 142128 800 142248 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 114006 180414 114062 181214 6 la_data_out[117]
port 262 nsew signal output
rlabel metal3 s 178270 154368 179070 154488 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 86314 180414 86370 181214 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal3 s 178270 129208 179070 129328 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 80518 180414 80574 181214 6 la_data_out[123]
port 269 nsew signal output
rlabel metal3 s 178270 159128 179070 159248 6 la_data_out[124]
port 270 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 la_data_out[125]
port 271 nsew signal output
rlabel metal3 s 178270 65288 179070 65408 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 66350 180414 66406 181214 6 la_data_out[12]
port 274 nsew signal output
rlabel metal3 s 178270 63928 179070 64048 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 170034 180414 170090 181214 6 la_data_out[14]
port 276 nsew signal output
rlabel metal3 s 178270 170688 179070 170808 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 72146 180414 72202 181214 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal3 s 178270 59848 179070 59968 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 62486 180414 62542 181214 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 156510 180414 156566 181214 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal3 s 178270 130568 179070 130688 6 la_data_out[23]
port 286 nsew signal output
rlabel metal3 s 178270 38768 179070 38888 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal3 s 178270 68688 179070 68808 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 100482 0 100538 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 157798 180414 157854 181214 6 la_data_out[29]
port 292 nsew signal output
rlabel metal3 s 0 128528 800 128648 6 la_data_out[2]
port 293 nsew signal output
rlabel metal3 s 178270 31288 179070 31408 6 la_data_out[30]
port 294 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 27066 180414 27122 181214 6 la_data_out[33]
port 297 nsew signal output
rlabel metal3 s 178270 91128 179070 91248 6 la_data_out[34]
port 298 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 la_data_out[35]
port 299 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 la_data_out[36]
port 300 nsew signal output
rlabel metal3 s 0 159808 800 159928 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 5814 180414 5870 181214 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 la_data_out[41]
port 306 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 la_data_out[42]
port 307 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 la_data_out[43]
port 308 nsew signal output
rlabel metal3 s 0 147568 800 147688 6 la_data_out[44]
port 309 nsew signal output
rlabel metal3 s 178270 37408 179070 37528 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 87602 180414 87658 181214 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal3 s 178270 71408 179070 71528 6 la_data_out[49]
port 314 nsew signal output
rlabel metal3 s 178270 146888 179070 147008 6 la_data_out[4]
port 315 nsew signal output
rlabel metal3 s 178270 166608 179070 166728 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 152002 180414 152058 181214 6 la_data_out[51]
port 317 nsew signal output
rlabel metal3 s 178270 145528 179070 145648 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 95974 180414 96030 181214 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 170678 0 170734 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 la_data_out[56]
port 322 nsew signal output
rlabel metal3 s 178270 78888 179070 79008 6 la_data_out[57]
port 323 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 la_data_out[58]
port 324 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 la_data_out[59]
port 325 nsew signal output
rlabel metal3 s 178270 117648 179070 117768 6 la_data_out[5]
port 326 nsew signal output
rlabel metal3 s 178270 96568 179070 96688 6 la_data_out[60]
port 327 nsew signal output
rlabel metal3 s 178270 165248 179070 165368 6 la_data_out[61]
port 328 nsew signal output
rlabel metal3 s 178270 135328 179070 135448 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 150070 0 150126 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal3 s 178270 138048 179070 138168 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 48318 180414 48374 181214 6 la_data_out[66]
port 333 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 43166 0 43222 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal3 s 178270 34688 179070 34808 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 43810 180414 43866 181214 6 la_data_out[70]
port 338 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 17406 180414 17462 181214 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 91466 180414 91522 181214 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal3 s 0 20408 800 20528 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 172610 0 172666 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 81806 180414 81862 181214 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal3 s 178270 121728 179070 121848 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 153290 180414 153346 181214 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 143630 180414 143686 181214 6 la_data_out[80]
port 349 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 la_data_out[81]
port 350 nsew signal output
rlabel metal3 s 178270 179528 179070 179648 6 la_data_out[82]
port 351 nsew signal output
rlabel metal3 s 178270 178168 179070 178288 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 125598 180414 125654 181214 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 9034 180414 9090 181214 6 la_data_out[88]
port 357 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 la_data_out[89]
port 358 nsew signal output
rlabel metal3 s 178270 19728 179070 19848 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 139122 180414 139178 181214 6 la_data_out[90]
port 360 nsew signal output
rlabel metal3 s 178270 36048 179070 36168 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 28354 180414 28410 181214 6 la_data_out[92]
port 362 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 la_data_out[93]
port 363 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 118514 180414 118570 181214 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 la_data_out[98]
port 368 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 la_data_out[99]
port 369 nsew signal output
rlabel metal3 s 0 171368 800 171488 6 la_data_out[9]
port 370 nsew signal output
rlabel metal3 s 178270 144168 179070 144288 6 la_oenb[0]
port 371 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 la_oenb[100]
port 372 nsew signal input
rlabel metal2 s 24490 180414 24546 181214 6 la_oenb[101]
port 373 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 la_oenb[102]
port 374 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 la_oenb[103]
port 375 nsew signal input
rlabel metal2 s 93398 180414 93454 181214 6 la_oenb[104]
port 376 nsew signal input
rlabel metal3 s 178270 111528 179070 111648 6 la_oenb[105]
port 377 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[106]
port 378 nsew signal input
rlabel metal2 s 132682 180414 132738 181214 6 la_oenb[107]
port 379 nsew signal input
rlabel metal3 s 178270 28568 179070 28688 6 la_oenb[108]
port 380 nsew signal input
rlabel metal2 s 79230 180414 79286 181214 6 la_oenb[109]
port 381 nsew signal input
rlabel metal2 s 173898 0 173954 800 6 la_oenb[10]
port 382 nsew signal input
rlabel metal2 s 12898 180414 12954 181214 6 la_oenb[110]
port 383 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 la_oenb[111]
port 384 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 la_oenb[112]
port 385 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_oenb[113]
port 386 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 la_oenb[114]
port 387 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[115]
port 388 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 la_oenb[116]
port 389 nsew signal input
rlabel metal2 s 25778 180414 25834 181214 6 la_oenb[117]
port 390 nsew signal input
rlabel metal2 s 130750 180414 130806 181214 6 la_oenb[118]
port 391 nsew signal input
rlabel metal3 s 178270 157768 179070 157888 6 la_oenb[119]
port 392 nsew signal input
rlabel metal2 s 18694 180414 18750 181214 6 la_oenb[11]
port 393 nsew signal input
rlabel metal2 s 35438 180414 35494 181214 6 la_oenb[120]
port 394 nsew signal input
rlabel metal3 s 178270 42168 179070 42288 6 la_oenb[121]
port 395 nsew signal input
rlabel metal2 s 7746 180414 7802 181214 6 la_oenb[122]
port 396 nsew signal input
rlabel metal3 s 178270 74808 179070 74928 6 la_oenb[123]
port 397 nsew signal input
rlabel metal3 s 0 136008 800 136128 6 la_oenb[124]
port 398 nsew signal input
rlabel metal2 s 57978 180414 58034 181214 6 la_oenb[125]
port 399 nsew signal input
rlabel metal3 s 0 167288 800 167408 6 la_oenb[126]
port 400 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 la_oenb[127]
port 401 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 la_oenb[12]
port 402 nsew signal input
rlabel metal3 s 178270 148928 179070 149048 6 la_oenb[13]
port 403 nsew signal input
rlabel metal3 s 178270 136688 179070 136808 6 la_oenb[14]
port 404 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 la_oenb[15]
port 405 nsew signal input
rlabel metal3 s 178270 123088 179070 123208 6 la_oenb[16]
port 406 nsew signal input
rlabel metal3 s 178270 67328 179070 67448 6 la_oenb[17]
port 407 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[18]
port 408 nsew signal input
rlabel metal2 s 97262 180414 97318 181214 6 la_oenb[19]
port 409 nsew signal input
rlabel metal2 s 149426 180414 149482 181214 6 la_oenb[1]
port 410 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 la_oenb[20]
port 411 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_oenb[21]
port 412 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_oenb[22]
port 413 nsew signal input
rlabel metal2 s 1950 180414 2006 181214 6 la_oenb[23]
port 414 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_oenb[24]
port 415 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_oenb[25]
port 416 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_oenb[26]
port 417 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 la_oenb[27]
port 418 nsew signal input
rlabel metal2 s 171966 180414 172022 181214 6 la_oenb[28]
port 419 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 la_oenb[29]
port 420 nsew signal input
rlabel metal2 s 126886 180414 126942 181214 6 la_oenb[2]
port 421 nsew signal input
rlabel metal3 s 178270 85008 179070 85128 6 la_oenb[30]
port 422 nsew signal input
rlabel metal2 s 141698 0 141754 800 6 la_oenb[31]
port 423 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 la_oenb[32]
port 424 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_oenb[33]
port 425 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[34]
port 426 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 la_oenb[35]
port 427 nsew signal input
rlabel metal3 s 178270 3408 179070 3528 6 la_oenb[36]
port 428 nsew signal input
rlabel metal3 s 178270 55088 179070 55208 6 la_oenb[37]
port 429 nsew signal input
rlabel metal2 s 42522 180414 42578 181214 6 la_oenb[38]
port 430 nsew signal input
rlabel metal3 s 178270 169328 179070 169448 6 la_oenb[39]
port 431 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 la_oenb[3]
port 432 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 la_oenb[40]
port 433 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 la_oenb[41]
port 434 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 la_oenb[42]
port 435 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 la_oenb[43]
port 436 nsew signal input
rlabel metal3 s 178270 101328 179070 101448 6 la_oenb[44]
port 437 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_oenb[45]
port 438 nsew signal input
rlabel metal2 s 111430 180414 111486 181214 6 la_oenb[46]
port 439 nsew signal input
rlabel metal2 s 154578 180414 154634 181214 6 la_oenb[47]
port 440 nsew signal input
rlabel metal3 s 0 178848 800 178968 6 la_oenb[48]
port 441 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_oenb[49]
port 442 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 la_oenb[4]
port 443 nsew signal input
rlabel metal2 s 160374 180414 160430 181214 6 la_oenb[50]
port 444 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 la_oenb[51]
port 445 nsew signal input
rlabel metal3 s 178270 150288 179070 150408 6 la_oenb[52]
port 446 nsew signal input
rlabel metal3 s 178270 62568 179070 62688 6 la_oenb[53]
port 447 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_oenb[54]
port 448 nsew signal input
rlabel metal2 s 141054 180414 141110 181214 6 la_oenb[55]
port 449 nsew signal input
rlabel metal2 s 34150 180414 34206 181214 6 la_oenb[56]
port 450 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[57]
port 451 nsew signal input
rlabel metal3 s 178270 116288 179070 116408 6 la_oenb[58]
port 452 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_oenb[59]
port 453 nsew signal input
rlabel metal3 s 178270 56448 179070 56568 6 la_oenb[5]
port 454 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_oenb[60]
port 455 nsew signal input
rlabel metal3 s 178270 7488 179070 7608 6 la_oenb[61]
port 456 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 la_oenb[62]
port 457 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 la_oenb[63]
port 458 nsew signal input
rlabel metal3 s 178270 81608 179070 81728 6 la_oenb[64]
port 459 nsew signal input
rlabel metal2 s 135258 180414 135314 181214 6 la_oenb[65]
port 460 nsew signal input
rlabel metal3 s 178270 167968 179070 168088 6 la_oenb[66]
port 461 nsew signal input
rlabel metal3 s 178270 9528 179070 9648 6 la_oenb[67]
port 462 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 la_oenb[68]
port 463 nsew signal input
rlabel metal3 s 178270 107448 179070 107568 6 la_oenb[69]
port 464 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 la_oenb[6]
port 465 nsew signal input
rlabel metal3 s 178270 172048 179070 172168 6 la_oenb[70]
port 466 nsew signal input
rlabel metal2 s 129462 180414 129518 181214 6 la_oenb[71]
port 467 nsew signal input
rlabel metal3 s 178270 21088 179070 21208 6 la_oenb[72]
port 468 nsew signal input
rlabel metal2 s 123666 180414 123722 181214 6 la_oenb[73]
port 469 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[74]
port 470 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_oenb[75]
port 471 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 la_oenb[76]
port 472 nsew signal input
rlabel metal2 s 18 0 74 800 6 la_oenb[77]
port 473 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[78]
port 474 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 la_oenb[79]
port 475 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 la_oenb[7]
port 476 nsew signal input
rlabel metal2 s 47030 180414 47086 181214 6 la_oenb[80]
port 477 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_oenb[81]
port 478 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 la_oenb[82]
port 479 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 la_oenb[83]
port 480 nsew signal input
rlabel metal2 s 90178 180414 90234 181214 6 la_oenb[84]
port 481 nsew signal input
rlabel metal2 s 50894 180414 50950 181214 6 la_oenb[85]
port 482 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[86]
port 483 nsew signal input
rlabel metal2 s 122378 180414 122434 181214 6 la_oenb[87]
port 484 nsew signal input
rlabel metal3 s 178270 48968 179070 49088 6 la_oenb[88]
port 485 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 la_oenb[89]
port 486 nsew signal input
rlabel metal3 s 178270 141448 179070 141568 6 la_oenb[8]
port 487 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 la_oenb[90]
port 488 nsew signal input
rlabel metal2 s 66994 0 67050 800 6 la_oenb[91]
port 489 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[92]
port 490 nsew signal input
rlabel metal3 s 178270 133968 179070 134088 6 la_oenb[93]
port 491 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_oenb[94]
port 492 nsew signal input
rlabel metal2 s 117226 180414 117282 181214 6 la_oenb[95]
port 493 nsew signal input
rlabel metal2 s 115294 180414 115350 181214 6 la_oenb[96]
port 494 nsew signal input
rlabel metal3 s 0 170008 800 170128 6 la_oenb[97]
port 495 nsew signal input
rlabel metal2 s 19982 180414 20038 181214 6 la_oenb[98]
port 496 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 la_oenb[99]
port 497 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_oenb[9]
port 498 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 user_clock2
port 499 nsew signal input
rlabel metal4 s 4208 2128 4528 179024 6 vccd1
port 500 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 179024 6 vccd1
port 500 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 179024 6 vccd1
port 500 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 179024 6 vccd1
port 500 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 179024 6 vccd1
port 500 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 179024 6 vccd1
port 500 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 179024 6 vssd1
port 501 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 179024 6 vssd1
port 501 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 179024 6 vssd1
port 501 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 179024 6 vssd1
port 501 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 179024 6 vssd1
port 501 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 179024 6 vssd1
port 501 nsew ground bidirectional
rlabel metal3 s 178270 87728 179070 87848 6 wb_clk_i
port 502 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 179070 181214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 48232444
string GDS_FILE /home/farhad/bin/Caravel_user_project/caravel_user_project/openlane/projtes/runs/22_09_10_23_16/results/signoff/projtes.magic.gds
string GDS_START 1105822
<< end >>

