VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO projtes
  CLASS BLOCK ;
  FOREIGN projtes ;
  ORIGIN 0.000 0.000 ;
  SIZE 895.350 BY 906.070 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 380.840 895.350 381.440 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 902.070 344.910 906.070 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 902.070 740.970 906.070 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 418.240 895.350 418.840 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 663.040 895.350 663.640 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 0.000 847.230 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 217.640 895.350 218.240 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.530 0.000 811.810 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 902.070 599.290 906.070 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 902.070 683.010 906.070 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 902.070 550.990 906.070 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 902.070 206.450 906.070 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 10.240 895.350 10.840 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 902.070 164.590 906.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 877.240 895.350 877.840 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 469.240 895.350 469.840 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 902.070 51.890 906.070 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 792.240 4.000 792.840 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 785.440 4.000 786.040 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 902.070 528.450 906.070 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 387.640 895.350 388.240 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 166.640 895.350 167.240 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 401.240 895.350 401.840 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.850 902.070 831.130 906.070 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 261.840 895.350 262.440 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 54.440 895.350 55.040 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 902.070 116.290 906.070 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 625.640 895.350 626.240 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.040 4.000 867.640 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 902.070 267.630 906.070 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 902.070 731.310 906.070 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 363.840 895.350 364.440 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 136.040 895.350 136.640 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.030 902.070 892.310 906.070 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 489.640 895.350 490.240 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.240 4.000 724.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 476.040 895.350 476.640 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 0.000 615.390 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 902.070 872.990 906.070 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 902.070 106.630 906.070 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 902.070 795.710 906.070 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 902.070 444.730 906.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 74.840 895.350 75.440 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 119.040 895.350 119.640 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 306.040 895.350 306.640 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 902.070 16.470 906.070 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 231.240 895.350 231.840 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 112.240 895.350 112.840 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 902.070 711.990 906.070 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 902.070 71.210 906.070 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 819.440 4.000 820.040 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 902.070 605.730 906.070 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 23.840 895.350 24.440 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 887.440 4.000 888.040 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 902.070 354.570 906.070 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 902.070 885.870 906.070 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 902.070 248.310 906.070 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 902.070 515.570 906.070 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 902.070 183.910 906.070 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 238.040 895.350 238.640 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 595.040 895.350 595.640 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 68.040 895.350 68.640 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 902.070 190.350 906.070 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 816.040 895.350 816.640 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 200.640 895.350 201.240 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 527.040 895.350 527.640 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 902.070 373.890 906.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 149.640 895.350 150.240 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 714.040 895.350 714.640 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 758.240 895.350 758.840 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.840 4.000 874.440 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 829.640 4.000 830.240 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 462.440 895.350 463.040 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 802.440 895.350 803.040 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 0.000 840.790 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.850 902.070 509.130 906.070 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 902.070 534.890 906.070 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 632.440 895.350 633.040 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 880.640 4.000 881.240 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 902.070 148.490 906.070 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 639.240 895.350 639.840 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 902.070 261.190 906.070 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 902.070 641.150 906.070 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 499.840 895.350 500.440 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 902.070 724.870 906.070 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 513.440 895.350 514.040 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 902.070 493.030 906.070 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 544.040 895.350 544.640 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 902.070 670.130 906.070 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 902.070 3.590 906.070 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 91.840 895.350 92.440 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 697.040 895.350 697.640 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.040 4.000 561.640 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 292.440 895.350 293.040 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 748.040 4.000 748.640 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 778.640 895.350 779.240 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 350.240 895.350 350.840 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 902.070 80.870 906.070 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 809.240 895.350 809.840 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 85.040 895.350 85.640 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 902.070 225.770 906.070 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 61.240 895.350 61.840 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 431.840 895.350 432.440 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 584.840 4.000 585.440 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 902.070 58.330 906.070 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 902.070 296.610 906.070 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 902.070 277.290 906.070 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 445.440 895.350 446.040 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 564.440 895.350 565.040 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 129.240 895.350 129.840 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 30.640 895.350 31.240 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 902.070 879.430 906.070 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 902.070 818.250 906.070 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 520.240 895.350 520.840 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.770 0.000 786.050 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 902.070 563.870 906.070 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 571.240 895.350 571.840 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 902.070 367.450 906.070 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 902.070 389.990 906.070 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 902.070 22.910 906.070 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.410 902.070 824.690 906.070 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 902.070 325.590 906.070 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 884.040 895.350 884.640 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 902.070 422.190 906.070 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 902.070 522.010 906.070 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 902.070 283.730 906.070 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 902.070 541.330 906.070 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.290 902.070 837.570 906.070 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.040 4.000 901.640 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 902.070 415.750 906.070 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 902.070 338.470 906.070 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 754.840 4.000 755.440 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 902.070 866.550 906.070 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 870.440 895.350 871.040 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 902.070 808.590 906.070 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 902.070 200.010 906.070 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 224.440 895.350 225.040 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 0.000 882.650 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 902.070 380.330 906.070 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 902.070 499.470 906.070 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 902.070 473.710 906.070 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 902.070 753.850 906.070 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 268.640 895.350 269.240 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 0.000 364.230 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 3.440 895.350 4.040 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 902.070 319.150 906.070 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 902.070 158.150 906.070 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 550.840 895.350 551.440 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 255.040 895.350 255.640 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 812.640 4.000 813.240 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 902.070 844.010 906.070 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 902.070 689.450 906.070 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 765.040 895.350 765.640 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 902.070 303.050 906.070 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 601.840 895.350 602.440 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 902.070 570.310 906.070 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 771.840 895.350 772.440 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 902.070 431.850 906.070 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 646.040 895.350 646.640 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 902.070 402.870 906.070 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 795.640 895.350 796.240 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 326.440 895.350 327.040 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 902.070 332.030 906.070 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 319.640 895.350 320.240 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 902.070 850.450 906.070 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 853.440 895.350 854.040 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 902.070 361.010 906.070 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 299.240 895.350 299.840 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 902.070 312.710 906.070 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 902.070 782.830 906.070 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 652.840 895.350 653.440 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 193.840 895.350 194.440 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 343.440 895.350 344.040 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 902.070 789.270 906.070 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 156.440 895.350 157.040 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 902.070 135.610 906.070 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 455.640 895.350 456.240 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 799.040 4.000 799.640 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 902.070 29.350 906.070 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 187.040 895.350 187.640 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 0.000 554.210 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 902.070 438.290 906.070 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 357.040 895.350 357.640 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 734.440 895.350 735.040 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 833.040 895.350 833.640 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 902.070 760.290 906.070 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 727.640 895.350 728.240 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 902.070 480.150 906.070 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 394.440 895.350 395.040 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 588.240 895.350 588.840 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 482.840 895.350 483.440 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 826.240 895.350 826.840 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 676.640 895.350 677.240 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 690.240 895.350 690.840 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.370 0.000 721.650 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 902.070 241.870 906.070 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 173.440 895.350 174.040 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 902.070 219.330 906.070 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 902.070 87.310 906.070 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 902.070 457.610 906.070 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 0.000 863.330 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 902.070 409.310 906.070 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 608.640 895.350 609.240 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 902.070 766.730 906.070 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 902.070 718.430 906.070 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 897.640 895.350 898.240 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 890.840 895.350 891.440 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 902.070 628.270 906.070 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 902.070 45.450 906.070 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 98.640 895.350 99.240 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 902.070 695.890 906.070 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 180.240 895.350 180.840 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 902.070 142.050 906.070 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 902.070 592.850 906.070 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 856.840 4.000 857.440 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 720.840 895.350 721.440 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 902.070 122.730 906.070 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.240 4.000 843.840 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 902.070 467.270 906.070 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 557.640 895.350 558.240 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 902.070 663.690 906.070 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 142.840 895.350 143.440 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 902.070 396.430 906.070 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 902.070 64.770 906.070 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 717.440 4.000 718.040 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 902.070 129.170 906.070 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 902.070 654.030 906.070 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 788.840 895.350 789.440 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 902.070 93.750 906.070 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 902.070 177.470 906.070 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 210.840 895.350 211.440 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 902.070 39.010 906.070 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 374.040 895.350 374.640 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 902.070 290.170 906.070 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 666.440 4.000 667.040 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 744.640 895.350 745.240 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 683.440 895.350 684.040 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 615.440 895.350 616.040 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 336.640 895.350 337.240 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 902.070 486.590 906.070 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 902.070 747.410 906.070 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 902.070 10.030 906.070 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 902.070 860.110 906.070 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 902.070 634.710 906.070 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 425.040 895.350 425.640 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 17.040 895.350 17.640 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 275.440 895.350 276.040 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 902.070 212.890 906.070 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 846.640 895.350 847.240 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 659.640 4.000 660.240 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 506.640 895.350 507.240 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 902.070 557.430 906.070 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 902.070 773.170 906.070 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 894.240 4.000 894.840 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 902.070 802.150 906.070 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 751.440 895.350 752.040 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 312.840 895.350 313.440 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 902.070 705.550 906.070 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 902.070 171.030 906.070 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 581.440 895.350 582.040 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 282.240 895.350 282.840 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 37.440 895.350 38.040 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 408.040 895.350 408.640 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 902.070 676.570 906.070 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 839.840 895.350 840.440 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 47.640 895.350 48.240 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 537.240 895.350 537.840 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 860.240 895.350 860.840 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 902.070 647.590 906.070 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 105.440 895.350 106.040 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 902.070 618.610 906.070 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 0.000 602.510 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.790 0.000 596.070 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 0.000 702.330 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 768.440 4.000 769.040 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 902.070 235.430 906.070 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 902.070 451.170 906.070 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.470 902.070 254.750 906.070 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.890 902.070 612.170 906.070 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 244.840 895.350 245.440 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 707.240 895.350 707.840 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 669.840 895.350 670.440 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 902.070 586.410 906.070 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 902.070 576.750 906.070 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 850.040 4.000 850.640 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 902.070 100.190 906.070 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 761.640 4.000 762.240 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 895.120 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 895.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 895.120 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 891.350 438.640 895.350 439.240 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 889.640 894.965 ;
      LAYER met1 ;
        RECT 5.520 8.540 891.870 895.120 ;
      LAYER met2 ;
        RECT 6.540 901.790 9.470 902.770 ;
        RECT 10.310 901.790 15.910 902.770 ;
        RECT 16.750 901.790 22.350 902.770 ;
        RECT 23.190 901.790 28.790 902.770 ;
        RECT 29.630 901.790 38.450 902.770 ;
        RECT 39.290 901.790 44.890 902.770 ;
        RECT 45.730 901.790 51.330 902.770 ;
        RECT 52.170 901.790 57.770 902.770 ;
        RECT 58.610 901.790 64.210 902.770 ;
        RECT 65.050 901.790 70.650 902.770 ;
        RECT 71.490 901.790 80.310 902.770 ;
        RECT 81.150 901.790 86.750 902.770 ;
        RECT 87.590 901.790 93.190 902.770 ;
        RECT 94.030 901.790 99.630 902.770 ;
        RECT 100.470 901.790 106.070 902.770 ;
        RECT 106.910 901.790 115.730 902.770 ;
        RECT 116.570 901.790 122.170 902.770 ;
        RECT 123.010 901.790 128.610 902.770 ;
        RECT 129.450 901.790 135.050 902.770 ;
        RECT 135.890 901.790 141.490 902.770 ;
        RECT 142.330 901.790 147.930 902.770 ;
        RECT 148.770 901.790 157.590 902.770 ;
        RECT 158.430 901.790 164.030 902.770 ;
        RECT 164.870 901.790 170.470 902.770 ;
        RECT 171.310 901.790 176.910 902.770 ;
        RECT 177.750 901.790 183.350 902.770 ;
        RECT 184.190 901.790 189.790 902.770 ;
        RECT 190.630 901.790 199.450 902.770 ;
        RECT 200.290 901.790 205.890 902.770 ;
        RECT 206.730 901.790 212.330 902.770 ;
        RECT 213.170 901.790 218.770 902.770 ;
        RECT 219.610 901.790 225.210 902.770 ;
        RECT 226.050 901.790 234.870 902.770 ;
        RECT 235.710 901.790 241.310 902.770 ;
        RECT 242.150 901.790 247.750 902.770 ;
        RECT 248.590 901.790 254.190 902.770 ;
        RECT 255.030 901.790 260.630 902.770 ;
        RECT 261.470 901.790 267.070 902.770 ;
        RECT 267.910 901.790 276.730 902.770 ;
        RECT 277.570 901.790 283.170 902.770 ;
        RECT 284.010 901.790 289.610 902.770 ;
        RECT 290.450 901.790 296.050 902.770 ;
        RECT 296.890 901.790 302.490 902.770 ;
        RECT 303.330 901.790 312.150 902.770 ;
        RECT 312.990 901.790 318.590 902.770 ;
        RECT 319.430 901.790 325.030 902.770 ;
        RECT 325.870 901.790 331.470 902.770 ;
        RECT 332.310 901.790 337.910 902.770 ;
        RECT 338.750 901.790 344.350 902.770 ;
        RECT 345.190 901.790 354.010 902.770 ;
        RECT 354.850 901.790 360.450 902.770 ;
        RECT 361.290 901.790 366.890 902.770 ;
        RECT 367.730 901.790 373.330 902.770 ;
        RECT 374.170 901.790 379.770 902.770 ;
        RECT 380.610 901.790 389.430 902.770 ;
        RECT 390.270 901.790 395.870 902.770 ;
        RECT 396.710 901.790 402.310 902.770 ;
        RECT 403.150 901.790 408.750 902.770 ;
        RECT 409.590 901.790 415.190 902.770 ;
        RECT 416.030 901.790 421.630 902.770 ;
        RECT 422.470 901.790 431.290 902.770 ;
        RECT 432.130 901.790 437.730 902.770 ;
        RECT 438.570 901.790 444.170 902.770 ;
        RECT 445.010 901.790 450.610 902.770 ;
        RECT 451.450 901.790 457.050 902.770 ;
        RECT 457.890 901.790 466.710 902.770 ;
        RECT 467.550 901.790 473.150 902.770 ;
        RECT 473.990 901.790 479.590 902.770 ;
        RECT 480.430 901.790 486.030 902.770 ;
        RECT 486.870 901.790 492.470 902.770 ;
        RECT 493.310 901.790 498.910 902.770 ;
        RECT 499.750 901.790 508.570 902.770 ;
        RECT 509.410 901.790 515.010 902.770 ;
        RECT 515.850 901.790 521.450 902.770 ;
        RECT 522.290 901.790 527.890 902.770 ;
        RECT 528.730 901.790 534.330 902.770 ;
        RECT 535.170 901.790 540.770 902.770 ;
        RECT 541.610 901.790 550.430 902.770 ;
        RECT 551.270 901.790 556.870 902.770 ;
        RECT 557.710 901.790 563.310 902.770 ;
        RECT 564.150 901.790 569.750 902.770 ;
        RECT 570.590 901.790 576.190 902.770 ;
        RECT 577.030 901.790 585.850 902.770 ;
        RECT 586.690 901.790 592.290 902.770 ;
        RECT 593.130 901.790 598.730 902.770 ;
        RECT 599.570 901.790 605.170 902.770 ;
        RECT 606.010 901.790 611.610 902.770 ;
        RECT 612.450 901.790 618.050 902.770 ;
        RECT 618.890 901.790 627.710 902.770 ;
        RECT 628.550 901.790 634.150 902.770 ;
        RECT 634.990 901.790 640.590 902.770 ;
        RECT 641.430 901.790 647.030 902.770 ;
        RECT 647.870 901.790 653.470 902.770 ;
        RECT 654.310 901.790 663.130 902.770 ;
        RECT 663.970 901.790 669.570 902.770 ;
        RECT 670.410 901.790 676.010 902.770 ;
        RECT 676.850 901.790 682.450 902.770 ;
        RECT 683.290 901.790 688.890 902.770 ;
        RECT 689.730 901.790 695.330 902.770 ;
        RECT 696.170 901.790 704.990 902.770 ;
        RECT 705.830 901.790 711.430 902.770 ;
        RECT 712.270 901.790 717.870 902.770 ;
        RECT 718.710 901.790 724.310 902.770 ;
        RECT 725.150 901.790 730.750 902.770 ;
        RECT 731.590 901.790 740.410 902.770 ;
        RECT 741.250 901.790 746.850 902.770 ;
        RECT 747.690 901.790 753.290 902.770 ;
        RECT 754.130 901.790 759.730 902.770 ;
        RECT 760.570 901.790 766.170 902.770 ;
        RECT 767.010 901.790 772.610 902.770 ;
        RECT 773.450 901.790 782.270 902.770 ;
        RECT 783.110 901.790 788.710 902.770 ;
        RECT 789.550 901.790 795.150 902.770 ;
        RECT 795.990 901.790 801.590 902.770 ;
        RECT 802.430 901.790 808.030 902.770 ;
        RECT 808.870 901.790 817.690 902.770 ;
        RECT 818.530 901.790 824.130 902.770 ;
        RECT 824.970 901.790 830.570 902.770 ;
        RECT 831.410 901.790 837.010 902.770 ;
        RECT 837.850 901.790 843.450 902.770 ;
        RECT 844.290 901.790 849.890 902.770 ;
        RECT 850.730 901.790 859.550 902.770 ;
        RECT 860.390 901.790 865.990 902.770 ;
        RECT 866.830 901.790 872.430 902.770 ;
        RECT 873.270 901.790 878.870 902.770 ;
        RECT 879.710 901.790 885.310 902.770 ;
        RECT 886.150 901.790 891.750 902.770 ;
        RECT 6.540 4.280 892.030 901.790 ;
        RECT 7.090 3.670 12.690 4.280 ;
        RECT 13.530 3.670 19.130 4.280 ;
        RECT 19.970 3.670 25.570 4.280 ;
        RECT 26.410 3.670 32.010 4.280 ;
        RECT 32.850 3.670 41.670 4.280 ;
        RECT 42.510 3.670 48.110 4.280 ;
        RECT 48.950 3.670 54.550 4.280 ;
        RECT 55.390 3.670 60.990 4.280 ;
        RECT 61.830 3.670 67.430 4.280 ;
        RECT 68.270 3.670 73.870 4.280 ;
        RECT 74.710 3.670 83.530 4.280 ;
        RECT 84.370 3.670 89.970 4.280 ;
        RECT 90.810 3.670 96.410 4.280 ;
        RECT 97.250 3.670 102.850 4.280 ;
        RECT 103.690 3.670 109.290 4.280 ;
        RECT 110.130 3.670 118.950 4.280 ;
        RECT 119.790 3.670 125.390 4.280 ;
        RECT 126.230 3.670 131.830 4.280 ;
        RECT 132.670 3.670 138.270 4.280 ;
        RECT 139.110 3.670 144.710 4.280 ;
        RECT 145.550 3.670 151.150 4.280 ;
        RECT 151.990 3.670 160.810 4.280 ;
        RECT 161.650 3.670 167.250 4.280 ;
        RECT 168.090 3.670 173.690 4.280 ;
        RECT 174.530 3.670 180.130 4.280 ;
        RECT 180.970 3.670 186.570 4.280 ;
        RECT 187.410 3.670 196.230 4.280 ;
        RECT 197.070 3.670 202.670 4.280 ;
        RECT 203.510 3.670 209.110 4.280 ;
        RECT 209.950 3.670 215.550 4.280 ;
        RECT 216.390 3.670 221.990 4.280 ;
        RECT 222.830 3.670 228.430 4.280 ;
        RECT 229.270 3.670 238.090 4.280 ;
        RECT 238.930 3.670 244.530 4.280 ;
        RECT 245.370 3.670 250.970 4.280 ;
        RECT 251.810 3.670 257.410 4.280 ;
        RECT 258.250 3.670 263.850 4.280 ;
        RECT 264.690 3.670 273.510 4.280 ;
        RECT 274.350 3.670 279.950 4.280 ;
        RECT 280.790 3.670 286.390 4.280 ;
        RECT 287.230 3.670 292.830 4.280 ;
        RECT 293.670 3.670 299.270 4.280 ;
        RECT 300.110 3.670 305.710 4.280 ;
        RECT 306.550 3.670 315.370 4.280 ;
        RECT 316.210 3.670 321.810 4.280 ;
        RECT 322.650 3.670 328.250 4.280 ;
        RECT 329.090 3.670 334.690 4.280 ;
        RECT 335.530 3.670 341.130 4.280 ;
        RECT 341.970 3.670 350.790 4.280 ;
        RECT 351.630 3.670 357.230 4.280 ;
        RECT 358.070 3.670 363.670 4.280 ;
        RECT 364.510 3.670 370.110 4.280 ;
        RECT 370.950 3.670 376.550 4.280 ;
        RECT 377.390 3.670 382.990 4.280 ;
        RECT 383.830 3.670 392.650 4.280 ;
        RECT 393.490 3.670 399.090 4.280 ;
        RECT 399.930 3.670 405.530 4.280 ;
        RECT 406.370 3.670 411.970 4.280 ;
        RECT 412.810 3.670 418.410 4.280 ;
        RECT 419.250 3.670 424.850 4.280 ;
        RECT 425.690 3.670 434.510 4.280 ;
        RECT 435.350 3.670 440.950 4.280 ;
        RECT 441.790 3.670 447.390 4.280 ;
        RECT 448.230 3.670 453.830 4.280 ;
        RECT 454.670 3.670 460.270 4.280 ;
        RECT 461.110 3.670 469.930 4.280 ;
        RECT 470.770 3.670 476.370 4.280 ;
        RECT 477.210 3.670 482.810 4.280 ;
        RECT 483.650 3.670 489.250 4.280 ;
        RECT 490.090 3.670 495.690 4.280 ;
        RECT 496.530 3.670 502.130 4.280 ;
        RECT 502.970 3.670 511.790 4.280 ;
        RECT 512.630 3.670 518.230 4.280 ;
        RECT 519.070 3.670 524.670 4.280 ;
        RECT 525.510 3.670 531.110 4.280 ;
        RECT 531.950 3.670 537.550 4.280 ;
        RECT 538.390 3.670 547.210 4.280 ;
        RECT 548.050 3.670 553.650 4.280 ;
        RECT 554.490 3.670 560.090 4.280 ;
        RECT 560.930 3.670 566.530 4.280 ;
        RECT 567.370 3.670 572.970 4.280 ;
        RECT 573.810 3.670 579.410 4.280 ;
        RECT 580.250 3.670 589.070 4.280 ;
        RECT 589.910 3.670 595.510 4.280 ;
        RECT 596.350 3.670 601.950 4.280 ;
        RECT 602.790 3.670 608.390 4.280 ;
        RECT 609.230 3.670 614.830 4.280 ;
        RECT 615.670 3.670 624.490 4.280 ;
        RECT 625.330 3.670 630.930 4.280 ;
        RECT 631.770 3.670 637.370 4.280 ;
        RECT 638.210 3.670 643.810 4.280 ;
        RECT 644.650 3.670 650.250 4.280 ;
        RECT 651.090 3.670 656.690 4.280 ;
        RECT 657.530 3.670 666.350 4.280 ;
        RECT 667.190 3.670 672.790 4.280 ;
        RECT 673.630 3.670 679.230 4.280 ;
        RECT 680.070 3.670 685.670 4.280 ;
        RECT 686.510 3.670 692.110 4.280 ;
        RECT 692.950 3.670 701.770 4.280 ;
        RECT 702.610 3.670 708.210 4.280 ;
        RECT 709.050 3.670 714.650 4.280 ;
        RECT 715.490 3.670 721.090 4.280 ;
        RECT 721.930 3.670 727.530 4.280 ;
        RECT 728.370 3.670 733.970 4.280 ;
        RECT 734.810 3.670 743.630 4.280 ;
        RECT 744.470 3.670 750.070 4.280 ;
        RECT 750.910 3.670 756.510 4.280 ;
        RECT 757.350 3.670 762.950 4.280 ;
        RECT 763.790 3.670 769.390 4.280 ;
        RECT 770.230 3.670 775.830 4.280 ;
        RECT 776.670 3.670 785.490 4.280 ;
        RECT 786.330 3.670 791.930 4.280 ;
        RECT 792.770 3.670 798.370 4.280 ;
        RECT 799.210 3.670 804.810 4.280 ;
        RECT 805.650 3.670 811.250 4.280 ;
        RECT 812.090 3.670 820.910 4.280 ;
        RECT 821.750 3.670 827.350 4.280 ;
        RECT 828.190 3.670 833.790 4.280 ;
        RECT 834.630 3.670 840.230 4.280 ;
        RECT 841.070 3.670 846.670 4.280 ;
        RECT 847.510 3.670 853.110 4.280 ;
        RECT 853.950 3.670 862.770 4.280 ;
        RECT 863.610 3.670 869.210 4.280 ;
        RECT 870.050 3.670 875.650 4.280 ;
        RECT 876.490 3.670 882.090 4.280 ;
        RECT 882.930 3.670 888.530 4.280 ;
        RECT 889.370 3.670 892.030 4.280 ;
      LAYER met3 ;
        RECT 4.000 897.240 890.950 898.105 ;
        RECT 4.000 895.240 891.350 897.240 ;
        RECT 4.400 893.840 891.350 895.240 ;
        RECT 4.000 891.840 891.350 893.840 ;
        RECT 4.000 890.440 890.950 891.840 ;
        RECT 4.000 888.440 891.350 890.440 ;
        RECT 4.400 887.040 891.350 888.440 ;
        RECT 4.000 885.040 891.350 887.040 ;
        RECT 4.000 883.640 890.950 885.040 ;
        RECT 4.000 881.640 891.350 883.640 ;
        RECT 4.400 880.240 891.350 881.640 ;
        RECT 4.000 878.240 891.350 880.240 ;
        RECT 4.000 876.840 890.950 878.240 ;
        RECT 4.000 874.840 891.350 876.840 ;
        RECT 4.400 873.440 891.350 874.840 ;
        RECT 4.000 871.440 891.350 873.440 ;
        RECT 4.000 870.040 890.950 871.440 ;
        RECT 4.000 868.040 891.350 870.040 ;
        RECT 4.400 866.640 891.350 868.040 ;
        RECT 4.000 861.240 891.350 866.640 ;
        RECT 4.000 859.840 890.950 861.240 ;
        RECT 4.000 857.840 891.350 859.840 ;
        RECT 4.400 856.440 891.350 857.840 ;
        RECT 4.000 854.440 891.350 856.440 ;
        RECT 4.000 853.040 890.950 854.440 ;
        RECT 4.000 851.040 891.350 853.040 ;
        RECT 4.400 849.640 891.350 851.040 ;
        RECT 4.000 847.640 891.350 849.640 ;
        RECT 4.000 846.240 890.950 847.640 ;
        RECT 4.000 844.240 891.350 846.240 ;
        RECT 4.400 842.840 891.350 844.240 ;
        RECT 4.000 840.840 891.350 842.840 ;
        RECT 4.000 839.440 890.950 840.840 ;
        RECT 4.000 837.440 891.350 839.440 ;
        RECT 4.400 836.040 891.350 837.440 ;
        RECT 4.000 834.040 891.350 836.040 ;
        RECT 4.000 832.640 890.950 834.040 ;
        RECT 4.000 830.640 891.350 832.640 ;
        RECT 4.400 829.240 891.350 830.640 ;
        RECT 4.000 827.240 891.350 829.240 ;
        RECT 4.000 825.840 890.950 827.240 ;
        RECT 4.000 820.440 891.350 825.840 ;
        RECT 4.400 819.040 891.350 820.440 ;
        RECT 4.000 817.040 891.350 819.040 ;
        RECT 4.000 815.640 890.950 817.040 ;
        RECT 4.000 813.640 891.350 815.640 ;
        RECT 4.400 812.240 891.350 813.640 ;
        RECT 4.000 810.240 891.350 812.240 ;
        RECT 4.000 808.840 890.950 810.240 ;
        RECT 4.000 806.840 891.350 808.840 ;
        RECT 4.400 805.440 891.350 806.840 ;
        RECT 4.000 803.440 891.350 805.440 ;
        RECT 4.000 802.040 890.950 803.440 ;
        RECT 4.000 800.040 891.350 802.040 ;
        RECT 4.400 798.640 891.350 800.040 ;
        RECT 4.000 796.640 891.350 798.640 ;
        RECT 4.000 795.240 890.950 796.640 ;
        RECT 4.000 793.240 891.350 795.240 ;
        RECT 4.400 791.840 891.350 793.240 ;
        RECT 4.000 789.840 891.350 791.840 ;
        RECT 4.000 788.440 890.950 789.840 ;
        RECT 4.000 786.440 891.350 788.440 ;
        RECT 4.400 785.040 891.350 786.440 ;
        RECT 4.000 779.640 891.350 785.040 ;
        RECT 4.000 778.240 890.950 779.640 ;
        RECT 4.000 776.240 891.350 778.240 ;
        RECT 4.400 774.840 891.350 776.240 ;
        RECT 4.000 772.840 891.350 774.840 ;
        RECT 4.000 771.440 890.950 772.840 ;
        RECT 4.000 769.440 891.350 771.440 ;
        RECT 4.400 768.040 891.350 769.440 ;
        RECT 4.000 766.040 891.350 768.040 ;
        RECT 4.000 764.640 890.950 766.040 ;
        RECT 4.000 762.640 891.350 764.640 ;
        RECT 4.400 761.240 891.350 762.640 ;
        RECT 4.000 759.240 891.350 761.240 ;
        RECT 4.000 757.840 890.950 759.240 ;
        RECT 4.000 755.840 891.350 757.840 ;
        RECT 4.400 754.440 891.350 755.840 ;
        RECT 4.000 752.440 891.350 754.440 ;
        RECT 4.000 751.040 890.950 752.440 ;
        RECT 4.000 749.040 891.350 751.040 ;
        RECT 4.400 747.640 891.350 749.040 ;
        RECT 4.000 745.640 891.350 747.640 ;
        RECT 4.000 744.240 890.950 745.640 ;
        RECT 4.000 738.840 891.350 744.240 ;
        RECT 4.400 737.440 891.350 738.840 ;
        RECT 4.000 735.440 891.350 737.440 ;
        RECT 4.000 734.040 890.950 735.440 ;
        RECT 4.000 732.040 891.350 734.040 ;
        RECT 4.400 730.640 891.350 732.040 ;
        RECT 4.000 728.640 891.350 730.640 ;
        RECT 4.000 727.240 890.950 728.640 ;
        RECT 4.000 725.240 891.350 727.240 ;
        RECT 4.400 723.840 891.350 725.240 ;
        RECT 4.000 721.840 891.350 723.840 ;
        RECT 4.000 720.440 890.950 721.840 ;
        RECT 4.000 718.440 891.350 720.440 ;
        RECT 4.400 717.040 891.350 718.440 ;
        RECT 4.000 715.040 891.350 717.040 ;
        RECT 4.000 713.640 890.950 715.040 ;
        RECT 4.000 711.640 891.350 713.640 ;
        RECT 4.400 710.240 891.350 711.640 ;
        RECT 4.000 708.240 891.350 710.240 ;
        RECT 4.000 706.840 890.950 708.240 ;
        RECT 4.000 704.840 891.350 706.840 ;
        RECT 4.400 703.440 891.350 704.840 ;
        RECT 4.000 698.040 891.350 703.440 ;
        RECT 4.000 696.640 890.950 698.040 ;
        RECT 4.000 694.640 891.350 696.640 ;
        RECT 4.400 693.240 891.350 694.640 ;
        RECT 4.000 691.240 891.350 693.240 ;
        RECT 4.000 689.840 890.950 691.240 ;
        RECT 4.000 687.840 891.350 689.840 ;
        RECT 4.400 686.440 891.350 687.840 ;
        RECT 4.000 684.440 891.350 686.440 ;
        RECT 4.000 683.040 890.950 684.440 ;
        RECT 4.000 681.040 891.350 683.040 ;
        RECT 4.400 679.640 891.350 681.040 ;
        RECT 4.000 677.640 891.350 679.640 ;
        RECT 4.000 676.240 890.950 677.640 ;
        RECT 4.000 674.240 891.350 676.240 ;
        RECT 4.400 672.840 891.350 674.240 ;
        RECT 4.000 670.840 891.350 672.840 ;
        RECT 4.000 669.440 890.950 670.840 ;
        RECT 4.000 667.440 891.350 669.440 ;
        RECT 4.400 666.040 891.350 667.440 ;
        RECT 4.000 664.040 891.350 666.040 ;
        RECT 4.000 662.640 890.950 664.040 ;
        RECT 4.000 660.640 891.350 662.640 ;
        RECT 4.400 659.240 891.350 660.640 ;
        RECT 4.000 653.840 891.350 659.240 ;
        RECT 4.000 652.440 890.950 653.840 ;
        RECT 4.000 650.440 891.350 652.440 ;
        RECT 4.400 649.040 891.350 650.440 ;
        RECT 4.000 647.040 891.350 649.040 ;
        RECT 4.000 645.640 890.950 647.040 ;
        RECT 4.000 643.640 891.350 645.640 ;
        RECT 4.400 642.240 891.350 643.640 ;
        RECT 4.000 640.240 891.350 642.240 ;
        RECT 4.000 638.840 890.950 640.240 ;
        RECT 4.000 636.840 891.350 638.840 ;
        RECT 4.400 635.440 891.350 636.840 ;
        RECT 4.000 633.440 891.350 635.440 ;
        RECT 4.000 632.040 890.950 633.440 ;
        RECT 4.000 630.040 891.350 632.040 ;
        RECT 4.400 628.640 891.350 630.040 ;
        RECT 4.000 626.640 891.350 628.640 ;
        RECT 4.000 625.240 890.950 626.640 ;
        RECT 4.000 623.240 891.350 625.240 ;
        RECT 4.400 621.840 891.350 623.240 ;
        RECT 4.000 616.440 891.350 621.840 ;
        RECT 4.000 615.040 890.950 616.440 ;
        RECT 4.000 613.040 891.350 615.040 ;
        RECT 4.400 611.640 891.350 613.040 ;
        RECT 4.000 609.640 891.350 611.640 ;
        RECT 4.000 608.240 890.950 609.640 ;
        RECT 4.000 606.240 891.350 608.240 ;
        RECT 4.400 604.840 891.350 606.240 ;
        RECT 4.000 602.840 891.350 604.840 ;
        RECT 4.000 601.440 890.950 602.840 ;
        RECT 4.000 599.440 891.350 601.440 ;
        RECT 4.400 598.040 891.350 599.440 ;
        RECT 4.000 596.040 891.350 598.040 ;
        RECT 4.000 594.640 890.950 596.040 ;
        RECT 4.000 592.640 891.350 594.640 ;
        RECT 4.400 591.240 891.350 592.640 ;
        RECT 4.000 589.240 891.350 591.240 ;
        RECT 4.000 587.840 890.950 589.240 ;
        RECT 4.000 585.840 891.350 587.840 ;
        RECT 4.400 584.440 891.350 585.840 ;
        RECT 4.000 582.440 891.350 584.440 ;
        RECT 4.000 581.040 890.950 582.440 ;
        RECT 4.000 579.040 891.350 581.040 ;
        RECT 4.400 577.640 891.350 579.040 ;
        RECT 4.000 572.240 891.350 577.640 ;
        RECT 4.000 570.840 890.950 572.240 ;
        RECT 4.000 568.840 891.350 570.840 ;
        RECT 4.400 567.440 891.350 568.840 ;
        RECT 4.000 565.440 891.350 567.440 ;
        RECT 4.000 564.040 890.950 565.440 ;
        RECT 4.000 562.040 891.350 564.040 ;
        RECT 4.400 560.640 891.350 562.040 ;
        RECT 4.000 558.640 891.350 560.640 ;
        RECT 4.000 557.240 890.950 558.640 ;
        RECT 4.000 555.240 891.350 557.240 ;
        RECT 4.400 553.840 891.350 555.240 ;
        RECT 4.000 551.840 891.350 553.840 ;
        RECT 4.000 550.440 890.950 551.840 ;
        RECT 4.000 548.440 891.350 550.440 ;
        RECT 4.400 547.040 891.350 548.440 ;
        RECT 4.000 545.040 891.350 547.040 ;
        RECT 4.000 543.640 890.950 545.040 ;
        RECT 4.000 541.640 891.350 543.640 ;
        RECT 4.400 540.240 891.350 541.640 ;
        RECT 4.000 538.240 891.350 540.240 ;
        RECT 4.000 536.840 890.950 538.240 ;
        RECT 4.000 531.440 891.350 536.840 ;
        RECT 4.400 530.040 891.350 531.440 ;
        RECT 4.000 528.040 891.350 530.040 ;
        RECT 4.000 526.640 890.950 528.040 ;
        RECT 4.000 524.640 891.350 526.640 ;
        RECT 4.400 523.240 891.350 524.640 ;
        RECT 4.000 521.240 891.350 523.240 ;
        RECT 4.000 519.840 890.950 521.240 ;
        RECT 4.000 517.840 891.350 519.840 ;
        RECT 4.400 516.440 891.350 517.840 ;
        RECT 4.000 514.440 891.350 516.440 ;
        RECT 4.000 513.040 890.950 514.440 ;
        RECT 4.000 511.040 891.350 513.040 ;
        RECT 4.400 509.640 891.350 511.040 ;
        RECT 4.000 507.640 891.350 509.640 ;
        RECT 4.000 506.240 890.950 507.640 ;
        RECT 4.000 504.240 891.350 506.240 ;
        RECT 4.400 502.840 891.350 504.240 ;
        RECT 4.000 500.840 891.350 502.840 ;
        RECT 4.000 499.440 890.950 500.840 ;
        RECT 4.000 497.440 891.350 499.440 ;
        RECT 4.400 496.040 891.350 497.440 ;
        RECT 4.000 490.640 891.350 496.040 ;
        RECT 4.000 489.240 890.950 490.640 ;
        RECT 4.000 487.240 891.350 489.240 ;
        RECT 4.400 485.840 891.350 487.240 ;
        RECT 4.000 483.840 891.350 485.840 ;
        RECT 4.000 482.440 890.950 483.840 ;
        RECT 4.000 480.440 891.350 482.440 ;
        RECT 4.400 479.040 891.350 480.440 ;
        RECT 4.000 477.040 891.350 479.040 ;
        RECT 4.000 475.640 890.950 477.040 ;
        RECT 4.000 473.640 891.350 475.640 ;
        RECT 4.400 472.240 891.350 473.640 ;
        RECT 4.000 470.240 891.350 472.240 ;
        RECT 4.000 468.840 890.950 470.240 ;
        RECT 4.000 466.840 891.350 468.840 ;
        RECT 4.400 465.440 891.350 466.840 ;
        RECT 4.000 463.440 891.350 465.440 ;
        RECT 4.000 462.040 890.950 463.440 ;
        RECT 4.000 460.040 891.350 462.040 ;
        RECT 4.400 458.640 891.350 460.040 ;
        RECT 4.000 456.640 891.350 458.640 ;
        RECT 4.000 455.240 890.950 456.640 ;
        RECT 4.000 449.840 891.350 455.240 ;
        RECT 4.400 448.440 891.350 449.840 ;
        RECT 4.000 446.440 891.350 448.440 ;
        RECT 4.000 445.040 890.950 446.440 ;
        RECT 4.000 443.040 891.350 445.040 ;
        RECT 4.400 441.640 891.350 443.040 ;
        RECT 4.000 439.640 891.350 441.640 ;
        RECT 4.000 438.240 890.950 439.640 ;
        RECT 4.000 436.240 891.350 438.240 ;
        RECT 4.400 434.840 891.350 436.240 ;
        RECT 4.000 432.840 891.350 434.840 ;
        RECT 4.000 431.440 890.950 432.840 ;
        RECT 4.000 429.440 891.350 431.440 ;
        RECT 4.400 428.040 891.350 429.440 ;
        RECT 4.000 426.040 891.350 428.040 ;
        RECT 4.000 424.640 890.950 426.040 ;
        RECT 4.000 422.640 891.350 424.640 ;
        RECT 4.400 421.240 891.350 422.640 ;
        RECT 4.000 419.240 891.350 421.240 ;
        RECT 4.000 417.840 890.950 419.240 ;
        RECT 4.000 415.840 891.350 417.840 ;
        RECT 4.400 414.440 891.350 415.840 ;
        RECT 4.000 409.040 891.350 414.440 ;
        RECT 4.000 407.640 890.950 409.040 ;
        RECT 4.000 405.640 891.350 407.640 ;
        RECT 4.400 404.240 891.350 405.640 ;
        RECT 4.000 402.240 891.350 404.240 ;
        RECT 4.000 400.840 890.950 402.240 ;
        RECT 4.000 398.840 891.350 400.840 ;
        RECT 4.400 397.440 891.350 398.840 ;
        RECT 4.000 395.440 891.350 397.440 ;
        RECT 4.000 394.040 890.950 395.440 ;
        RECT 4.000 392.040 891.350 394.040 ;
        RECT 4.400 390.640 891.350 392.040 ;
        RECT 4.000 388.640 891.350 390.640 ;
        RECT 4.000 387.240 890.950 388.640 ;
        RECT 4.000 385.240 891.350 387.240 ;
        RECT 4.400 383.840 891.350 385.240 ;
        RECT 4.000 381.840 891.350 383.840 ;
        RECT 4.000 380.440 890.950 381.840 ;
        RECT 4.000 378.440 891.350 380.440 ;
        RECT 4.400 377.040 891.350 378.440 ;
        RECT 4.000 375.040 891.350 377.040 ;
        RECT 4.000 373.640 890.950 375.040 ;
        RECT 4.000 368.240 891.350 373.640 ;
        RECT 4.400 366.840 891.350 368.240 ;
        RECT 4.000 364.840 891.350 366.840 ;
        RECT 4.000 363.440 890.950 364.840 ;
        RECT 4.000 361.440 891.350 363.440 ;
        RECT 4.400 360.040 891.350 361.440 ;
        RECT 4.000 358.040 891.350 360.040 ;
        RECT 4.000 356.640 890.950 358.040 ;
        RECT 4.000 354.640 891.350 356.640 ;
        RECT 4.400 353.240 891.350 354.640 ;
        RECT 4.000 351.240 891.350 353.240 ;
        RECT 4.000 349.840 890.950 351.240 ;
        RECT 4.000 347.840 891.350 349.840 ;
        RECT 4.400 346.440 891.350 347.840 ;
        RECT 4.000 344.440 891.350 346.440 ;
        RECT 4.000 343.040 890.950 344.440 ;
        RECT 4.000 341.040 891.350 343.040 ;
        RECT 4.400 339.640 891.350 341.040 ;
        RECT 4.000 337.640 891.350 339.640 ;
        RECT 4.000 336.240 890.950 337.640 ;
        RECT 4.000 334.240 891.350 336.240 ;
        RECT 4.400 332.840 891.350 334.240 ;
        RECT 4.000 327.440 891.350 332.840 ;
        RECT 4.000 326.040 890.950 327.440 ;
        RECT 4.000 324.040 891.350 326.040 ;
        RECT 4.400 322.640 891.350 324.040 ;
        RECT 4.000 320.640 891.350 322.640 ;
        RECT 4.000 319.240 890.950 320.640 ;
        RECT 4.000 317.240 891.350 319.240 ;
        RECT 4.400 315.840 891.350 317.240 ;
        RECT 4.000 313.840 891.350 315.840 ;
        RECT 4.000 312.440 890.950 313.840 ;
        RECT 4.000 310.440 891.350 312.440 ;
        RECT 4.400 309.040 891.350 310.440 ;
        RECT 4.000 307.040 891.350 309.040 ;
        RECT 4.000 305.640 890.950 307.040 ;
        RECT 4.000 303.640 891.350 305.640 ;
        RECT 4.400 302.240 891.350 303.640 ;
        RECT 4.000 300.240 891.350 302.240 ;
        RECT 4.000 298.840 890.950 300.240 ;
        RECT 4.000 296.840 891.350 298.840 ;
        RECT 4.400 295.440 891.350 296.840 ;
        RECT 4.000 293.440 891.350 295.440 ;
        RECT 4.000 292.040 890.950 293.440 ;
        RECT 4.000 290.040 891.350 292.040 ;
        RECT 4.400 288.640 891.350 290.040 ;
        RECT 4.000 283.240 891.350 288.640 ;
        RECT 4.000 281.840 890.950 283.240 ;
        RECT 4.000 279.840 891.350 281.840 ;
        RECT 4.400 278.440 891.350 279.840 ;
        RECT 4.000 276.440 891.350 278.440 ;
        RECT 4.000 275.040 890.950 276.440 ;
        RECT 4.000 273.040 891.350 275.040 ;
        RECT 4.400 271.640 891.350 273.040 ;
        RECT 4.000 269.640 891.350 271.640 ;
        RECT 4.000 268.240 890.950 269.640 ;
        RECT 4.000 266.240 891.350 268.240 ;
        RECT 4.400 264.840 891.350 266.240 ;
        RECT 4.000 262.840 891.350 264.840 ;
        RECT 4.000 261.440 890.950 262.840 ;
        RECT 4.000 259.440 891.350 261.440 ;
        RECT 4.400 258.040 891.350 259.440 ;
        RECT 4.000 256.040 891.350 258.040 ;
        RECT 4.000 254.640 890.950 256.040 ;
        RECT 4.000 252.640 891.350 254.640 ;
        RECT 4.400 251.240 891.350 252.640 ;
        RECT 4.000 245.840 891.350 251.240 ;
        RECT 4.000 244.440 890.950 245.840 ;
        RECT 4.000 242.440 891.350 244.440 ;
        RECT 4.400 241.040 891.350 242.440 ;
        RECT 4.000 239.040 891.350 241.040 ;
        RECT 4.000 237.640 890.950 239.040 ;
        RECT 4.000 235.640 891.350 237.640 ;
        RECT 4.400 234.240 891.350 235.640 ;
        RECT 4.000 232.240 891.350 234.240 ;
        RECT 4.000 230.840 890.950 232.240 ;
        RECT 4.000 228.840 891.350 230.840 ;
        RECT 4.400 227.440 891.350 228.840 ;
        RECT 4.000 225.440 891.350 227.440 ;
        RECT 4.000 224.040 890.950 225.440 ;
        RECT 4.000 222.040 891.350 224.040 ;
        RECT 4.400 220.640 891.350 222.040 ;
        RECT 4.000 218.640 891.350 220.640 ;
        RECT 4.000 217.240 890.950 218.640 ;
        RECT 4.000 215.240 891.350 217.240 ;
        RECT 4.400 213.840 891.350 215.240 ;
        RECT 4.000 211.840 891.350 213.840 ;
        RECT 4.000 210.440 890.950 211.840 ;
        RECT 4.000 208.440 891.350 210.440 ;
        RECT 4.400 207.040 891.350 208.440 ;
        RECT 4.000 201.640 891.350 207.040 ;
        RECT 4.000 200.240 890.950 201.640 ;
        RECT 4.000 198.240 891.350 200.240 ;
        RECT 4.400 196.840 891.350 198.240 ;
        RECT 4.000 194.840 891.350 196.840 ;
        RECT 4.000 193.440 890.950 194.840 ;
        RECT 4.000 191.440 891.350 193.440 ;
        RECT 4.400 190.040 891.350 191.440 ;
        RECT 4.000 188.040 891.350 190.040 ;
        RECT 4.000 186.640 890.950 188.040 ;
        RECT 4.000 184.640 891.350 186.640 ;
        RECT 4.400 183.240 891.350 184.640 ;
        RECT 4.000 181.240 891.350 183.240 ;
        RECT 4.000 179.840 890.950 181.240 ;
        RECT 4.000 177.840 891.350 179.840 ;
        RECT 4.400 176.440 891.350 177.840 ;
        RECT 4.000 174.440 891.350 176.440 ;
        RECT 4.000 173.040 890.950 174.440 ;
        RECT 4.000 171.040 891.350 173.040 ;
        RECT 4.400 169.640 891.350 171.040 ;
        RECT 4.000 167.640 891.350 169.640 ;
        RECT 4.000 166.240 890.950 167.640 ;
        RECT 4.000 160.840 891.350 166.240 ;
        RECT 4.400 159.440 891.350 160.840 ;
        RECT 4.000 157.440 891.350 159.440 ;
        RECT 4.000 156.040 890.950 157.440 ;
        RECT 4.000 154.040 891.350 156.040 ;
        RECT 4.400 152.640 891.350 154.040 ;
        RECT 4.000 150.640 891.350 152.640 ;
        RECT 4.000 149.240 890.950 150.640 ;
        RECT 4.000 147.240 891.350 149.240 ;
        RECT 4.400 145.840 891.350 147.240 ;
        RECT 4.000 143.840 891.350 145.840 ;
        RECT 4.000 142.440 890.950 143.840 ;
        RECT 4.000 140.440 891.350 142.440 ;
        RECT 4.400 139.040 891.350 140.440 ;
        RECT 4.000 137.040 891.350 139.040 ;
        RECT 4.000 135.640 890.950 137.040 ;
        RECT 4.000 133.640 891.350 135.640 ;
        RECT 4.400 132.240 891.350 133.640 ;
        RECT 4.000 130.240 891.350 132.240 ;
        RECT 4.000 128.840 890.950 130.240 ;
        RECT 4.000 126.840 891.350 128.840 ;
        RECT 4.400 125.440 891.350 126.840 ;
        RECT 4.000 120.040 891.350 125.440 ;
        RECT 4.000 118.640 890.950 120.040 ;
        RECT 4.000 116.640 891.350 118.640 ;
        RECT 4.400 115.240 891.350 116.640 ;
        RECT 4.000 113.240 891.350 115.240 ;
        RECT 4.000 111.840 890.950 113.240 ;
        RECT 4.000 109.840 891.350 111.840 ;
        RECT 4.400 108.440 891.350 109.840 ;
        RECT 4.000 106.440 891.350 108.440 ;
        RECT 4.000 105.040 890.950 106.440 ;
        RECT 4.000 103.040 891.350 105.040 ;
        RECT 4.400 101.640 891.350 103.040 ;
        RECT 4.000 99.640 891.350 101.640 ;
        RECT 4.000 98.240 890.950 99.640 ;
        RECT 4.000 96.240 891.350 98.240 ;
        RECT 4.400 94.840 891.350 96.240 ;
        RECT 4.000 92.840 891.350 94.840 ;
        RECT 4.000 91.440 890.950 92.840 ;
        RECT 4.000 89.440 891.350 91.440 ;
        RECT 4.400 88.040 891.350 89.440 ;
        RECT 4.000 86.040 891.350 88.040 ;
        RECT 4.000 84.640 890.950 86.040 ;
        RECT 4.000 79.240 891.350 84.640 ;
        RECT 4.400 77.840 891.350 79.240 ;
        RECT 4.000 75.840 891.350 77.840 ;
        RECT 4.000 74.440 890.950 75.840 ;
        RECT 4.000 72.440 891.350 74.440 ;
        RECT 4.400 71.040 891.350 72.440 ;
        RECT 4.000 69.040 891.350 71.040 ;
        RECT 4.000 67.640 890.950 69.040 ;
        RECT 4.000 65.640 891.350 67.640 ;
        RECT 4.400 64.240 891.350 65.640 ;
        RECT 4.000 62.240 891.350 64.240 ;
        RECT 4.000 60.840 890.950 62.240 ;
        RECT 4.000 58.840 891.350 60.840 ;
        RECT 4.400 57.440 891.350 58.840 ;
        RECT 4.000 55.440 891.350 57.440 ;
        RECT 4.000 54.040 890.950 55.440 ;
        RECT 4.000 52.040 891.350 54.040 ;
        RECT 4.400 50.640 891.350 52.040 ;
        RECT 4.000 48.640 891.350 50.640 ;
        RECT 4.000 47.240 890.950 48.640 ;
        RECT 4.000 45.240 891.350 47.240 ;
        RECT 4.400 43.840 891.350 45.240 ;
        RECT 4.000 38.440 891.350 43.840 ;
        RECT 4.000 37.040 890.950 38.440 ;
        RECT 4.000 35.040 891.350 37.040 ;
        RECT 4.400 33.640 891.350 35.040 ;
        RECT 4.000 31.640 891.350 33.640 ;
        RECT 4.000 30.240 890.950 31.640 ;
        RECT 4.000 28.240 891.350 30.240 ;
        RECT 4.400 26.840 891.350 28.240 ;
        RECT 4.000 24.840 891.350 26.840 ;
        RECT 4.000 23.440 890.950 24.840 ;
        RECT 4.000 21.440 891.350 23.440 ;
        RECT 4.400 20.040 891.350 21.440 ;
        RECT 4.000 18.040 891.350 20.040 ;
        RECT 4.000 16.640 890.950 18.040 ;
        RECT 4.000 14.640 891.350 16.640 ;
        RECT 4.400 13.240 891.350 14.640 ;
        RECT 4.000 11.240 891.350 13.240 ;
        RECT 4.000 9.840 890.950 11.240 ;
        RECT 4.000 7.840 891.350 9.840 ;
        RECT 4.400 6.975 891.350 7.840 ;
      LAYER met4 ;
        RECT 27.895 44.375 97.440 885.185 ;
        RECT 99.840 44.375 174.240 885.185 ;
        RECT 176.640 44.375 251.040 885.185 ;
        RECT 253.440 44.375 327.840 885.185 ;
        RECT 330.240 44.375 404.640 885.185 ;
        RECT 407.040 44.375 481.440 885.185 ;
        RECT 483.840 44.375 558.240 885.185 ;
        RECT 560.640 44.375 635.040 885.185 ;
        RECT 637.440 44.375 711.840 885.185 ;
        RECT 714.240 44.375 788.640 885.185 ;
        RECT 791.040 44.375 820.345 885.185 ;
  END
END projtes
END LIBRARY

